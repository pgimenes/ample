`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
I0n7NAh7lPD9ghjhTWY7q5FVi1iLeBFtNrwfbxJCCTGbv7hyrzRl82B5+WKGS0KB8dT7KOh5qgE2
LpTWFkOceg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fUGxIqWLpkp7p+hgpMfaT86uYBfXa6tnZz/bjWOgnj91tJIjZ4HMCD4MAtgfmK0x2Xpe5Wb7NLPO
s87MSCVVCBiOA/h3SGBbCl6+SJr8kvCbH5F9/bvYCmN4uXqxsxbhKq22KWEHZToxndnWcctbnRQn
35ocXUo0D1o26tLxWwU=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MiaF3K4Km1PZq1kKcMCaubE/GNIkpr17yqdcPEkVH/mWCIEANuarAwQyZdqvJorYhunwizVbbQFD
FjZP2gz8WOcBuMRfJrrCVkBMcbBKnquInJyzCj/0qVbPulJ1P30gFehdTHRWAp7lWhez5WUllMuk
kUnBmgLdkb/EuE+DmBm7tyUqExPjQbjgUljP1Ut6Yd6swb7QD1OEJ1wk0BEopAMOueco4FaEcRml
u+POHgZQALby1FcEK+8BR+tXtedWu0DLDAjLEiI2c8Kd4Us6zn29oaATqNYzanhrdYgTSOwM+PE3
Z+oqOVYKom9pea7iP67dNwTYsbLLWunrz5jsOg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
spgx6sVCkLoyQGrTVoM0LLggqZcOWIYUTQpk1U2Q7QSZUxoZSlAesqGt8a7ujG01ww9BGpt7ArAD
LVZh88WY1tAVX82jnKzh7QuPNMfNI4WwKVkJI3CiQzEusVBtQ4M1fPBKItUzEvyA0+QUtTXS5Rp5
G+LLF0CqHqlsxQBWxABQ0rpRc1NNrs8ktfDtO5o8pEDRUcG8mrdH6sSlqnk0PDzsti92TfgChXf9
+P/D7KzGFstMLoTdavEG+fHKAnHbeX/Yf4LGHm9pfqyNg2pTGnapfa8vm5o9UMVCzocco9WSvCsj
doa+2gFH2v1jFtXZgOh1Pfinpf6mNIVEvrTpmg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
l5uAZd91bKvtCPTGfKStVfJ/YcQwPEc1QJSpTy2G1IZaFGkZ2VuNDR6Wcj1roY27HhOWV8Yd1whL
/f9j1AntqRTxMpfOkX8XdZZOONq5w7+Mdp6O7eRbBunGuCfnuTq2ysecwCzdBvAWC3VI2NAs8lrX
3mNW74wwKWzhpShZv/1T1bC+8slNmlm8YHeC/5xvRaIPvXewkTQ5WWQEVQ/WSutnuy/3/ZQRbUSi
PSsS/KRuDp034MGeSvQcxDceYeyXqZjJFUua1j6rww+/8pglaSklFowRq29p24zU+8wjQjvRveC1
HkDsqQScm4Qv3f0xsoo/slaciZypQ+rDZ6TQXA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
c+DB3pUEAuBFXd1H3t+yms0J2EMKNwI3jBYkWMq+YxHY4XgO4QSU1vC1CpvU6oHyQk/h6yOgD5N+
V6eZb2aAuMa1b1aYdeeo5zHszJZWHWuSqw+qjw8iD2wuJ9lZ98W28ZVvHcbcJM2MZ89WJ2aKjKba
+WosNIUVJ1mNKhv7OVs=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WCYIyMJb9GXyx3NLwNdDRIsLlZMjmFag8BCvf+pcuxC4FtORBfd/r3l1IkUQR231iCqLPDCl5AMF
aJcZKwNHm0YYti1t4+5bKHmwQWRPa3J2D+yCVjH1cV1BuJazU/xZqaemQPB0dIgFfOP4ZkbttE5I
Tg5YEN4YAPMZAhZN6hyfTuWiU8749sHYa6d2Ox1iHm3B5GyU6HOXKXZWg+UgbtVT7rR5IQecGZHG
sbZ5DpjlPLob0w+ctwr/o8Kmn/Jo1zFIpCXnBIaVUVnyvAOGE63/K/W66tmOkSYxwF6GIUoZ6kVR
sPw4+MrbxZn/xPQh/DOGe2geS1PV/uZrzRQSSA==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
wISAlnbnTQHiY1JyL4+OR/F6r17CVXaNVzt1ojURbmsRII6P0rjnXmQi0pHB9nDaMakKiQIS/6jl
a/IM7qMNhC4rxshGk8FkR84FiTb5kaNXnxVRd+DjcQr6p2kyBXYea4u7oUQ5Wsa4AynUfNe6W+bP
Xe0mC8Dfpli5JCAIv6GTufCytdIF5p61TKUs8eP8pWlSq0U1tzrriS28H4Cu6W69UK8KQcKCRLr9
8Tk/ggkLrbs+bSuHBdv9hGyyNJi0WZZk8pk/8HpYFFoTNQkcfL8kSDRMNJvvQRmkc6UVwH3zeE3f
ki/RBQIhr7A7610ZCWRBAVGj2EHh7N4rKw4fvg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
EfreCivSIJjH8rlCp+zLAPX5molEG565xFicuIc9iMRik86yt/s44rc81so/RRm6h/FZDb4urn4m
YdT5jMEPhIU5Td7TXHIp6CR4hpH8sZLRSqP4nyfqGVBXl3PT3usY3IOoAxaZGCMWDlAHxqfZ5EXZ
AnzYxuOmyudAKPytymw5SqBEEewXCPmwVOOz0b301LSXtKIxnpvFVMpKw7J/9IOJlBhTY+mNRVqs
gu6h3xAVt61fLU7otYdQ7K+t3sKDttaJufqiwvR8EZDdPfKhdekoBK2kRJCzoJx/w74pFZ0OFI6n
fZEZIW8Zly5AWQ2Lx8xSDbyPhUAbLtoGjIOkHvNwNcdegq6WSsp/Ds34n9a6P4qg4d+M5JHjdWNy
ndd/Z1jnNEk97GpfqYezHO1TlizJO2juEoPtFNxfIR3gO6k3y6btuJiEWaSDhw0BfhR+pFiQP80k
hVv66hHpanBKFKdl5gkcniGU2zhZ4x+ObSbYsfFNgcCIiRZ0tkDwpcggowxVtQ9ctuGHUMzbUony
xq2m/qyFFo6YJlYRqWD258KuWTkjei1Dpyaegv9xiGYZ+FcY+DhmpbibBuToCWgSAxq6UWGv7Fcp
o2NxFnY/qpsZBSArodHenaYasc3/R3bRSnIvn9eLmUaa5ZRQoqKeHXY8QrUK/YcYKaQF2GhlAvus
iOAwZPW7YNSFaW1mIvW999POIT8rdokMZoK7LDJ70ptc/r543FSAoEjlptReoHcSpJwr0z1w/8YG
LpWM9tQEr8Syk/k36OLOK1cNQXWij7QvEWM9RBI/KPKR1v9art6WjaWPSMZGzyZxBSu6ZLHUQO3H
skXJ+SZknsd/KdX4PwIVR2MlVOyD/MuPHniP5gO5KqWtDomt4uLJgNMfbWekzVlEvMRJOKx5tpEe
cgrelQu3xp+HZ+8UcLcXAOnRGH1MB9dluXt1Tih+wULziL2OXlvTZUUBRZ48PEB/fW0sRUxOHr0O
xsdfFMN0ar6hAAlIr+CNrxggdH3kqJ2OvlC5hHcX1BoOPgz3Z1kq7rsp7Mf5OxfJnob5Vco8lW9S
IHDm1eJpD/0jhLyUHrvF7uWDlzD3dc3iPrw9oeLiv+drsfRHGpUilqlDk+F6Kq49FZTY3x86jUNE
ZS5FLNJTyIyiHSqxvR63Bh1Eb2Pb1NY6e54IY1e6JECyfGado9TL0XJxPsloUUnDtPxH4Lu2K0fa
ULr/JPP5XplEeFaf2rfQZhd7xvYivlez99T+raRyYH/oRgh6HgRPVQgHCE0OINSM/U+ebuSwtN9u
xUkt9AZ7B/UWs0NrqHehpsmp04yqUnQfpd4fU0b5FUK6S8s6dY2pW77yyrMGpEJdPZxVJOWkB/y+
TcuibamDenWWp7F3o+cNJ/Ronawk2szOmL2yObPylalZwvUYM8cZuRjyUyuUlA2/1mq9oWUvOeXS
8YbHkwanPiiOw2WGLrpTngsTgVRYmdlAyXTPfgOgtAn1d2PeK/RJBhDY0NlNGFy+3SaUKcyeYMBS
FWc+NB0v3RpGXXT0w+23L6tzD9As4UR5zRWV+hCuIPhZiCwEBHUVSNrNei06Nmbh/yw7HHRCtNr7
wFfcG1xdlcWYEizPsOX+NHi6eO+eisgW7CC6IrBlBV/qCRKnxNQUe06ydg+fEzysgQVgQw7xvI10
JElehrkpU27Yo3TcgZM3UILs7gwJoNznjy6KmnNEaUogxEpoD6E5nge8vDpztLg/cbO6PZQ8DYRU
ILQA93oUuE9dWGYFUr2xcCWIC4DZYdWJNqwe6ptwI9Hy/Q6GZyRphdVjRqSaBBjmIk1cev0qNTML
ypoNMOdZ3sn8XcdVIv8ZsBGCkZ7mZHAqh8QsT/VkkX4kSQuOz2+AijcH380fsxrM3QHTA+eN54Ez
h01qlPHQFhNA7qvDeBi8vWyq4jUuCDcx+tn/X2f2W8pBqfdsJU0faRedjlgWWN1wbglW1mRWOdT+
yqB42zlVnnY6XmxbWGgWVIbsX9wkpmCnFRwd363cXc5RLkMaYWqFO4+UfSOS/fklQuX7bBlzaZ1L
uBpqV1NBIGeR+d7Zsq0wfM4O0flPFdlCJoz5oRXFSoYhVdm28OVWtVn/fzOb50GSCBnsvpz2SkU3
NZAvgi74+UEiDT/V5GShAJOd+7OO8o2qHxhj0lkWInWG1RQW7UsErYM5YiEE2BX/pFXRoEAjaqNU
LYmDRZ3Oo0ATfRPTL9QDz+sn6rgOEoFDVCxoyO2TcTG6axxfni+4c4r0AAqPcWdMSR3yduMaImO1
SPU4Gcc/xn7kx1XBNdkU5M1Ql4NnT85pIL8YR3bwEK7hF6OU+QZBJKnzkys+W+WUaATW6spUJuCI
OZN4i4JE55D186B4Dn6a6I3Z1vxZw3538SHSGcBcpkZU0d+XfTPgeSFHOVlwKcKqEJo76wyft7wd
4gnPY/CiJ35gA2nirpo2kymPxLhWtsYFx1giRYwb5uKxWbt5Fl+FgeBzm1gFHEH1oG5D09X9e9rT
KUSuQ5J2AjTklbgQwh9InxpcnDw5cwrBiBdukGI0xqRNKNyMSPs85cmIgyty3meEOPUbVL4X9KFZ
nPgyBGzET0qAeoV0lVQejQVpUreUL78gQYEF7XU7UmpQQHV7qzUAMazs4PpxXjBY2PRyFuqc6pmP
8PIMAp2vpTH6wdX+GEj0BqqbhPT+cCL1ccUmsFd+bGrVciSfMcSuRDkgnXvF+szKe40rUSBcqJ6O
EUrKaW1scWLc7esjeZ5vsk0XQVaipzPev4Qb5pL+kV3fZl84Q4JmSiISflF07fk/lKAEfaboX+jF
hLcQG9Q5AAYyBLK4Dol/hnbERTYkgFooZ3QVZgXrO0fgNkoBXaZDzIm2TniKdlkOM+f3on1oBfjw
tjABcMAZasnJGoX3JGu78ijEizvs3OPCzZsfb8zwoj/cEz8r2i5nxZ08X9y3/GoTe1i3oWsJrnCL
YtNfp5bJTV5BDyAGICDQvq64FFh0Fd4MpGeTNLv/CVGAOV8m6rRIsiyKwXs6D+e14wiEKw+5PkRg
I4GSK3vvEXn+TCvpEz7JeySUipiuM7a//lQL0LevU583c55gpKGCpEJSHJz/sLDnZ/DSuLFs/mHI
Vm+c1cI2SXz8og69I79rFI2eg8NiysEAglcszXZR3TEC+XZ2q9h/Hfl/6KIbGQ6qFmirvtg/o5T1
Z2gIC2MyBGpKMD/n6mAw8P0Efz8aqptk473jP5FHsG1DYjCT7Vh6QGT05TU+QnynlJg6dZlvNB3e
y+Hdr+wMgaUBxSbRAhMNnjdpg6/vduIhS11DHu8DLCFzykbrDAbCYzfc3zMh7nE+H4G3WqI4ElDI
Ii+lUzEA5dFKx7k6hCNNAW7WyPl4EeEQtK9hi/+RT8HxBu7oON102MVgignDaCLE6jSasmVVgPUK
5RvQOpTMvhVNJ1O6+bpnbIl3RZnqeHOqbnpveQJZhrJGYMV1/WrdnFQayEGaH206Jx9qpSRQgf00
Y1cNEpc0lQzLPdL/2E1JlGAbNBji0uEKJBa8pYewQkj6Q4V3baxzXJo2pzcU5e0fpxOUl8qOUcVa
lbkaeMrBG2b441ZurX0GR2yopfpVyIUNF8Plp8qV8Kg1kjOYbpgPYGiPT7Oh75TRAbzKzkfSMuAh
sHWWZD6pwYrBzDysEsT58gl8iPgpSVCY1NpebvfwVnj0YHle8oaGmQ/C4vjs2gOTUHdsNz57H6Nv
s28oNS1cMh3/iUVJadZec5nEyKXu6frl84vb86i/QNbM7jqK3gOcFBWCSptAhiZXN1L8/Gc2l4Js
JSQNqEQJILpvUNy+K7PB79kiRGDSzBbZ2aXFoCVtQSq9Qymgl1EthiTqYTpznR4W9YqiPUzWyhjC
jZ2PxtijLh6cxGzWt1q2jOC/AU3GLqFv1A9em8fBnRxnPqa+zEPUNXgBtDNfRFcoZ9c9sKP0E47H
SSim65sQVUwGvjpurCH912HTsHYxL4gJgbCQcgXLiJLk1YybZbQI0PhrT2q7OjnP6EzVncBJ0QIB
HGWTce/xW/YSQtifBhcxfHF59s+O4k1buVWdBw/t2zvI/aayqWry1/ClkHqlj2lFpkW0Sxy1mbW+
YTNyrUlT3tytpMaFLF8qLZAwn1wJrKX/V4MFBNoqEIj7ri43/ntKjh2cPihPdbD5OJKuX5HsxcBn
sNshUbmpSJWpDiidvygkB+3K+x6EDzsE4GcamGENY2g2mw6+/Dd+XVj4PKylTWR5hEAIqnZHl9Ws
wcayOr26/caqPOyu5NwKjHh03TVzO0Y/JvUTaeGXvFgS034uJWLoZm2WFvNJI1qBRJ4Zg/5MOa7G
mKOu/30z98+7PQqc8krYtDh+0/Q9KHcVxr8qg3frGafSNOCoR3fKo4ltQb3SPorTwAatli82i2jI
r2ULPxS0vZWjqMm2Z/t5GJnVeGE6XnQoao3cnQaK5gHb8wb3EUSUBdhvSxB2vnVg1vY17WEMtBN1
KZWik0BJXCAnWgB/lYuYnSwGJsJgdyjPPabrlL2YiyX0kQrhsNZ4/ogN8+YiC5rRp9OGH7cMSG+s
fQ+EAHsqNCa0iRLEm/V23YJbSnxxHyk51047qlBtOao9dp+0vXHaDL70GVOKSSMie3TNrGWTGLx5
xCeFTsWQQOCY0YrFffLSCxBz6XTnlkxaKw09Lqq43c9j3Q+sWlf2qZ571grXDqILk2GcHhnD9hBZ
/hUsX6mKocl8yODHK9rMDV793mRLw0L68ByNtZnwupJvICAhdalrkGg4NSDnvZCuD4xVl/jsa0Q+
87WUFE3j4XdYjjLjFKAeYQEAKfu//5gVPPQPhHswFvGNQvU/3WtKqbsYtcW/IrWwGgZ0LxflljeU
3wnf6T+AJ8rvGkJpoK3zu2HrgcJtUDXsLuB8UthKUH9+cAGM/CRjv50WYFTZASR18YGrbEzfQW7d
HPhMW5Cm7470VA+D5LpL+N6O5lGcHFh6i84WQPInS9nCHFBH9nlC69HC8IZlfIb+nDBeqKQVAwZx
u1FiMhc7ewvGlItzMtJtSv2O8y87BjXBinLXvYd3f4CWYaVrLF/e1kpGFNTe9Jbt2PuuVggZIIJo
nAlgAk/ObSalfmfx0COh4OePF7ZQwt8MTqHWKXjumTwZcd3wQHuZmbbBO4egVaNosd/hmKbgSM5W
Mv1CNRWAKbjolAeAg/92khKGK0kT6gmgVdG+fzk3Y7IGOGpOs2canPSAXiKClQ1ZuBpaoalfA8td
sVnvCpCx6COnwEAL48fWC7q+YIEXMOjyR+2pYkdEHsZV7GqBDbktKW09RDiJNZiGx9+C8KJrpBGK
2oMycL4skePV3e2MLwuzs86YFVq4NFYel6sklCNVDJdnj96aqfPc6Ewhg8ncwJfXjhUEKEKxh8Xn
e9ownUkC9UOBe/x7tdMaRLFtqVQu+1hefISNSkfu0EXUS42cUNUom/pkOvRCh/OpBPq9A2G5weKa
/bfcE9EdRfZ/Ek1sFW8G7uaDIXD8W3SUVrXFXKwTkf35INitKL5KtLPLN9TN1zrj6Ok+tABjUEbB
3G1c+L/FpdtdRiE6Qc+Bkz8gvgQXGRHFepxIrpYjNK7v3yaLY7MtDSbyXyIJuixrDeRpqCn5LFkN
TrbKJDi38A6orS3FOjxjhdY3aw9R81xmJyX9A80/eZjfrL0RhCQFPCEoIthmy8LyVFYIN62xIjlx
ytUt6ypWpBg1Pr27gM2X7uQTqj6wej1w8AwAuYRVEo7Kv4C/6wzSi2HMmeC4rDlHjDZdiybQMSrZ
AIhjKuSvrvn6GUBoG6rAVabcoDCe9W/L6KGc5Um5W2X2KhF7XP8HC01FURDPI74DT0QAMNm5QBd3
pEETE3Hd1bfCk3xd5pdqJ2BXxrALH2raGuY8VNq4el5l3N0Es5Kmp/QIlKE80xu3XhSRnyoGiVOI
iwduYfooCXE8GsSEKToYR8A04wlQreQZZfuJKy2TxMP2GIJ+76j9vJbSW3zJUUKVlwT4XSYCCMqs
fxwrdoGyyroluqx8YQTkRn5RDlbPfi9MhFIqlqvIeMrCyjmqrf8aUeIGumskq6CaYZABez9oP/0i
CkliUNWSRLiorUQJCPWIAmT+pt4llClby4+0cB4awG2Eqqox0E9SEeE/JVGegHHwoJy2ujdSyKHn
oo30Vp9dtvjPZYIX/ad1QfpofM0V/p52qn9uAQFZbFXKROCtPUrekC64z5B1dAo1TQSVdeUnXcRs
KQytL7/rCmj0AVko/BcDGRGaA5/0ocNUWNGC1bnEdlo/34Q4RmZtWTic45WYb+GdowL24Pt20f6V
Ea1CnsoEY4sFN/ZgAJtEHK8GehmK0cyPKkjqFHaNMkoia7s8Ol4YNo28Om6euKuV2CtvCNjgMOJ2
tY433Z2WmPGd9yym7VbTQpcj7dhyaSvY0Pw1IDzs7sO4D4yXjGybiKXCNtrsE2Db3iC/hRtHzs8U
9M9cpG+tx704Myv9R2tFYHUtsI4B2mbBbQBTCftPYq1UwfuIsaMYQwr8JnYPmhrH3VspwbJUWK1p
j7h5bLwmExJLAiz5yI9C5kjf3LQ/IGowJr82AWyoKMe1IULun4bUnhMhq+JXE1RqH5sI6UHtxNcG
vB4ioYJLKbghngm//hk21HToCczAYOgwJkUd+uqPcp+eBi3KTm96p1EiNriEs1u+C5ydce1r1cM3
0Q4b9V57vlh7mHoFF0JfHgYE5PUqhPLOyEG1D4UMENluY9Cf7edywq2mDmK1xImXFOrTMzIqlzeD
1SUSrcc1TMsH2/Qmkg+KWO6OLbCkUd5PlWDA0XOlpLz5WiUG3r7xTfxMF2TLgbb8aSqDjpKyhxNa
+RsFeW4ErnfKgMBHXwh45+YLH+CaRh55qjYxosER4dCrI6ife6P1F2lwz6sdlMGuYW197fFVgnGk
8VSlHC5mfLPSvqQJQJRwNkQUdE7272WPl5uj5pJ7ec89lpatPYu8xf/a19ilaBJ4AM2jau/ziCn2
iSs+ZiVdPC5+kBtgYKfr6kylAfm1su7z26zUC+EcRPil9tGFBJQwdvFma30AhBy4QhrV5QpCpa57
6w2TW0++IytlM90W+uXAHjxMk/V5PlaQrfocx5xdV/ZWEekEIVcOQfOTwjC1zGTVth9g1IuV8INR
+LmUgRuVTKVpt0IXhzKYPBsdLaXeqAFSlSuJ9pwdzcAc7UqyVCr/K4if4expADlQkM08CniJxnpb
id0QAj6CIvEZfHx809IEvTdm0zdPYekOYdn+BLq+EEbEYD2MCyCHGTsojmkwEOZCkZ7IASsfvgBL
vd6EtTFKXu3MeG1cklAyLGpupXd/yTUDB1BCRTYW82NvC3ZGbEYRzMi7TVSkWxL/dbrrp3xnt0pR
hk9uPORO1c3LO0D7/VvpdmVHO1U4TRa4xSfHgzskNeKd/bqDqOxQcv57pVHPFvi3ToAdF14s12QH
KGZPFL42J6wSjzA/yL90fiobFJlupm2Rl1jYc6Y8BXbzGdGrZshbTbf/bwvcZfAeQpIoA4aHOG4w
+9SQU/Z+dTaI+OjrN9caeylprP8gOsoMh2LaiG7+b2g3Ul+1f+LNYcIJ4Sqd38PZ7AIysAG6RPZ8
JOh/+PiASQRI0/SgmuTsfhV7kgMHzNavXIpflt629kN+/9Ak+53BdRNjuuwIznJ3qBvmVfjz6taf
/paUnTwewLdPzTPMzTa60tGdRaRUqBmNiNg0LQkCrZcyzE62h/pCyxDZb/L+ErUnrQ0w2q43shxq
kKi5ww67l2L97+SRBSktoUmU9ITZLlRU/nrmGQ5OFfwVNMTTlvHWcOqJjfd3yEA3Tol8le79OTeo
VXwwwBzuSjNBBtYb2XleEDVnjHOXzoEVw88+pKwte9lqsLvBs+qrygh314iptxdHF4rJhPW0EK9R
lflAo4zE8WUPX9lQ8yJ3b72l00rdP6e4utlIQZN7JuANaMuABBK87we7+N0Jy+AJrBXPuwMOhRSj
QQEBlZXeZq7JkNsCdugCBAXlGqxLzFdlhVVMAhFWy6u8bNshP6XNZl8BwDU3TLffmei9M3dtT1HT
zRWbV/B0vgyVGr7rqX8E7cwdJq8X/XGU6mqcCkbCljoJEakCMllYrauzPLXla8Ex9ipV4drblG9q
9X2GHF0QSg4cFLywL3fvXx11etiAfRarWER3Dp632s+NwRX1cUbK/4R/ScllCEHDKQxrDCML+dMr
Z7ccyOPJpNiteknczb06GwAwzDXZCKlOQfew+oMs9yUDfMsPlPDmRmxzHIgX9tOP+tqaX8tUmBLn
gHEb9rqsVw2bROIOnWOnCEWttH6xY4d1I3gUBXQ8zcJ9QYGDPTjYv3jpMeT9FFPz4OtGsJF3M6di
LESAfcFVO7ZYQrMkX5lY2mIwpHUQ5n6fx39C5Tg3w6/am773kB8Ys+leL9f8YB8Dypgo86EiGMhu
ZaPon+m+fv1G1AJVDRsXxXrunDF0Ta0D1NXAGuxzyp6CnWrRkmQ1Cc78Q1r3WvErYe+uE5Kq5FAZ
gu7JvqmOla6OvIudDNmHkWm8g35lMAnAwS1tivjWgdYVipQluKENzPSRHllUCVL/dolzoSnVxjSe
cSWntn9JEGWov/q7jS6ugjt6ByuhQQAIHL7F3E+Dz8YGEVENidVXV5BDKLMzu0A/2HXeiHhdZHxy
YHcKVqaHcqZXFAoLOQMolVAC3gB7ygF7OlQQRZhHufzllfP1MfeMpqhBkT/kv/78Vx9bbyNyJMFB
vCgXojB78EwmE18FaRpO0km5DdUQdYJClbs/sOgAls2AZ6Fshh5E73JJ5167YLfJi0xE/Vk+BSAd
eL4P76QPfZgalDC4hEZmxZJOeTU/Qky+L4342lIqpb1GHk9AuDZCpFvV97JkESdBQeJkz+biZCji
IoN9KGywbbD5bKNSK4eTr3MBbtpnGqPkoeyJXhUglB7Ha4LUlyTyySfKodjyt5eAetGQNPiCO0Mk
W+yhSYMeGjWdZPg1ROfVSL2z9ikt1D7wAQlF18ol5tlL69K9HA3hTbwKQnHrbsQYpkj6Gf92IF+P
c34TaQYRZOo+WXKnh0Y7dU676rXLGg7Fzexb7FsI2c2JxN+V544X/sTsC6OkPgerlL5pndCfXtKv
0DtBpk5ia/Fi6lwSNb/2NQhGFemFnkLDtQHyKhXopCDf37Uy9LCCMlelpLMEGaz5EelOWJ0X/3p1
evJX/ia8FOzr1sIu5WHu+VOi7LQ56VWHXSqbsN5fUcNv033FiE+AYHkJte12ZHRfoVu/ccfvZnDc
tY9ZWiucY/JmYHtNVLrcQRZS/K5K0em/e8dnoa7XAQyKC7XixaPD2+tuDJWOf6OJAwdlkeNyAtrH
mn8xeUxRde8f7YFI1NPAus/hFvUjt0d/GNdAwMdiRRiq4EwCzzOBAvtp+1YzT2UEaAkTdfaTK467
QS/aTXWVEv5iKP8rQCgKvYZCAsU++XNZcEYrnDjm2m0YaahvhFikyFVH3F0EoQp0zYGlPoOHJ3cU
pSvy/kXDilJn6RnQ1aQhEBHKmXBT4/lNPPt6WFGkfBswvdRvqBvlWY8jezR9GCQt7IQ2yFNmjvZQ
mTMpwFQC1++41RyKk2r2hyuRRbuhGE4KjJvc/pZ6BWCN8W6j6fNlafusRbX5hquk7SEBGLNKyzX5
ROuPdSHOvy787sKUW46+R3ViHcv9BkhVyDJ8FN2ReJyusmlXAW2xDWyaKZ6o0PAvcidPDLRGh1FE
6gdGRoD3zfQKnhCmG/x5kYo+NsfT9dlN7FR3++ZygU6ET/lO2tBWoSk2zPTlcZ9f79+SGpElo1Rj
nBmRVM/gSVZq3rxjLS9/DZXSQ7b192JMrws4I2AffhTi+cjZD0DmgMb0T4MoFKq3QOQz1zVGn/u7
zF5zciJI4FBvUXzAXlSX4h/JKyGEtsNYcoe480oyZGiRmzu37A6c2bQC81fmuq5tI5wmXj0rmEMH
JqpH9IQFWy0dUoSu/K+efAFz+CuatbP3bvG+7ErjdzYDMR6R6LMvOMBpKHjse81vRAxN34vEiHVy
BoRr89h793TnjU2ungN6lrwnQ84B4V54s8fN4aAlsq3c/4DBdkiNFOvBBZ8/olGXuOJrisayMewk
TMf1CzhLeLb/G9KrIlp2f9VIKsFlcKDvTx0i0c4LztzQ54scagqi5+eT8Ypx2DD3c71NE71CkAjU
dYEkvxF2K86qsV+mZL5lbsRcOcJvsYME/Yqdo7SGKwt25XbzXN/e4ooDzv8CDpNSs/lOhqTmVO62
3Wo/CTN2ogJirJbHUwN1QpxCvmvKbn+k7XuY7gmpJNAOXLsIPdtriUr3nAFfufEqS4vT+1jQMOc3
pyRl6dTIXNJALO6HamRdIlw7GCmOke2gjMSE8ixZ+YSxEDyZ6CvMUx/oPi04rixjPFL/SZ26/72n
8wffsOpfhK58DPezCHrpSqNpQOQ/1uItV1sLIzyD2DMGeILIrFLAZSmE7n41EJMzla019v59UDoO
aLUF38kmqxs0cA2v9bOtRU+x56nnlNv0h6PIHyS4QRKwuMR/ptYvaIkqp8EHsPZP2H2e9zIbe33X
9RKVMR19UuzN40pqOpre19BwhZBL0HziyiwNRYO1ByvCA461xHHotDy4eMp4/0Ag0wcE02Otm46M
x9GwsGylQg2xBCxPQ+EP1UNosHTKWm8AyXOlqYQ2smLUYit903LwoTLY5AMOAT0+O+txD9qdSxv5
WJaAD43+TY1BdWaN+q6W7P+EhDDhH/Dfava6sYF7ZINX7dPRrFGK91TU28/ep3P3m7NOJ+7AOQ3Q
bWk4h9hYDNB0mRAssUefbEWuImfgtG3a/QgJfyYp0uRA8RiH5SpQG9nCTdi+fjGumPAWXiR4mL5y
yTyTVrdz8yY9JPWnsY/IYZAYIQT/jqOkQC0FALegAa0ShiYfqO4UyQqc+vInC4gmyaqUN40QX+Ig
TOXXtV2ef9SsD6qqDdYIfEHQj0Df828arglqV2Q7mOs6WOgB7xcEv4Wdm22OkZMCF5ob3YAUdWnG
DHJpQQ6uwEIYTOLjuHSuFQiWzlaqd5lBwJU+yVn4UKpVMSTkCGwPLXc+2dXman8l+n6ROTMaQ76o
EHro3NuVMM9slH4fUiZNHkIThJcaPQz/tWMfUsJ538CdjYaBWlGhDJ2rgc5k9PyBBT/nLYTqsI8h
ahgBhf+1J+0fnH+xAC+ddaORPuvrCKL3EtX2F/paf0amGvfDxpA61YQ0/PH9woeHtDKlkb02Ii/B
cx0tg4l4t4nc4cSsQpJpabt6u9as6zmohPfm02i+nYB/z9DnUj8T9q4sR3Mr3S/+IK4zFaCsDhTt
st9a9d0WvJ6tu0QVwNLZ8nWjSXmaKvWkLpmduUaqEuqCoubMZCqPRH+FtDq7zcT52sRspGUVqNq2
xGCNA/UkCtqclckbTuLMRbmX9cOvfIyasAZqrp0SwGstMWjPZm+JVHI1Sks74AXu+DY4lLYe/pij
T2N/NpQ8lwdD5J9KFrHH6I3q53hFze/DQBHRiEJrpVrHEQgR00sRQ1w+Gncuyv+KtsOYkw1GoMc5
Ghh4zDAaFRoZIEvPuu3qtJej2wCDM2Kz+HQyParRaPnCBdlcVGLvcPb9HsJgxBhXGlg1/sQ6NMKI
GIpEovQfCY/fgZsAqOkA4vAZaP6PNb00Ist0aurJP73IvtzzcmTxUnaTPxeyD+eN2y79/ws1ZXxm
u3/IRWTg7SED34ffRdgdIw7N5+R1FBGb3ec6loEijjFDh25gt5p8greE8VepXZlQ9WXfb7t6cbDn
4oVJyrpSWEmhUxfKPK2HYc18rRlbnL4iUh0JnIatO9vn5p86UgnpAvY0uh42QI3igxQ03eAT6bZz
bsv7cjCIrqp1F6XX4MAy9gn8nFWd01aeWUyEqsLinRzuul6+GpP8wP87bIeP4El/CPLxQ6166FZc
EjvJoKP3e8XJqCYDezr8CQiOweIu9o36BYkG/pKmWrD2yyZRe+Un7aLkDiWRsOSS9tzMPwVx9foV
YWBI8/BwQggJTP8uTew6WQ6HQxUzYuZCcFly17FVJjzMWt261kXuqFiylrqrGGKM+xNRiIfu62G4
p16xLad5eQ87vd4XoM/A4nC083bKhSD7yRs97vZ0rXxxhyJrGwP69mb7H1aXag3u3nLeTb2xgHhA
upvrkmmDJL8EE2tq+OcODbj8H1ez+xMFeue8+UJwqYKRrO2AqymBP4OxlnwdTJm2whz+sFesIh/N
PeaNFEo8L+p2zy/AR0Bwi3WIDlrONKwAQHp7GZTI9Pi/UpcpIQjhKMJ6WIRhgHAthMZk1mYTDfHa
1RMB4Zjr1ZK3mgQQpTE5gs7r2UgnQVrnagfFgB5vVtG3BC91kkKhiVlqjM7HzLX7wo5+YtWYob1P
bSjgKP3XegQeOcEKaI0BkR74oPiqxdHXvwOtgPCsVAW7QC5R+ydqmZ1tzp24phZIdT5cJerrp1RZ
NDT6NoJyCESNlYH2EAPn095GtLftJdtZtDT4LiBZmqPwsMPbo7hlFWEhE78YgvZtW9Pr2pq9XQSJ
cIF5EHpzjkz94HMPHUn9bkJcDcOVs5fs81i24b3udFVIGRdRnc0OyaKo03eWQY6fTXJV2J1xH1i7
fa3f4H4plcPGg752jwBV6aXqkJPZYKBLml427XLgewXNTHZnJ0rh+fSAIJpbcVWNKqRkInSNo5pU
l+RzJDDrDGEmC68SA2SwSiGjIPb1NS0xgH/EjOokBl1pWLzfnKnGefRDV398Hj9oAsllAxA0XZNQ
4/uYneZZ0IuYfDz7xI/ZMuYTbh4LW7CJgHd3xTcbCIle9LI30FNgM68HYV6a5eJj8foEu1gwp9Ng
Gf7fM270vGKDBnAspwTgnOEWCLYKG3pEK9hKU0l02v5ClJy7ReR7Wm5VCuxftCWi0stnyVkPB2zk
FScfehyP6Yf5cxmc9Z4M2tWC4gJ3Y8jHu6GM8UW5XH72Lafr56GOy8u05Y+Yv7ANK8UBltD2dR2J
CjKD1rB6nMD7rJk7BQjXViGX9+vJZrGALIToXArLFjrxgOJWitcZSxcmozHh2WtBZqHgLEBvsqTJ
hg1Om6hGO8F9hzBE3HkI4Wf9rlBAxWZKG6z8OSWy1jgvAWM7T29Q/DeHQR+gQ/IFDGjeyobbSJtk
3Q3AQPU8sDsh2AgUL0/jbMr395haKL3XSc2qkGtkfVfQ4j8HBlsIZ4y/tqv8YDvFqUgv8H0h9J7D
7x8hLzQFdNAVYHb7K13GniBxCFS4LzrsEoHgprLBlcrHunhDZCHKpeySC1Kdrz6hULIbT3pthRg+
6j0cqrYJPjTEQOQR7S88tggY2WrPGLSrM7xj659WbAvodUi1wK1wlCjBQ/RbLNkaSijpElxoCNVX
MI+d4MMnL1BFrkQs4AmYtlAe9t4ey+bPHyAsNpz9R78z4aPw5CUL2EDay+vqmqUAeNVELpCWwQrv
OpcP2YhaWGcebMODcLZ4dDHKiC2ltpTeKB+gwkqe27GpEQfL8qTkv/VicInk10ddGBmR7X0f1hTX
+0egboYpA+2QjsLQcCppsSRHyJG2G3Yn15Hmargs/oV16lVHX7PbrEGH4yxK3pKvuiCROII6tmY3
D/ycrXALthjvmA0QSOLLpjLbeHiNPng9OpSjJlI+8fUfi5DN2JlRsoS6f7gotwh2+Mnp9mjwq1gm
WlP5ye2oafCWrDxTOeaeSCiq1oI5pUhYg74jya1j9u+Mbkf8xM1ecDgmBSCgnduVm/oiHDH4Bf1C
5YYn1UD1qyGcobGj3PR08r+1XJEFi4Ug6n/Ftr+Mv/ahgQMbZnmcXI7vpaZM5mMGR+6ZnU917FFC
7g8mRh0kUeLLExm2jc7T2xyW69+NukboQ7WGVxZ77aSrq0CmF+IHy9UTMEAVPBL4iob9SJpbg3LO
lCIIkpdJ1G/GgEack4rMxSEd6JpiCN1hj7q9kFROjyIxHFT3j2H49o/rO8aDVNUQzBv+3ypWOKPP
Rd1682HwGTVfrKjJqoIpF+65yGHG5Mo4S5rCFAqZuTogFmlhNdzwVsrdmPpMGAXIkESEoaIkN0s4
s714EgQ8rLCzfiNQSgCAlWtc1aDaQJNtD21+Q0EH2PY4i3ODkgEpzFWjs5vTleXi6NCidsphbm36
HilzEYbqRPLoJqy3E1uWzd8svD7CnZli8I+xp4AGwsn93dSWKPfbKmVkcC/ogCsTdWH5Jdc9D9AK
c4qh0C8PQGQF0IfWjttDUMjdz7uW3E94iP9JUTlgwUBUP6cZlBroBxsDd+sisMLRrjIWvmm2gnL6
ZjVLiBJ43TcaNfRwZmIRM+JswonoSm1vE1LSFq3rhUY5syMaJVL4+sdMSPejhSisX4mPh7JTQKKZ
gGE0qNfKiC1I81QVcPaTN1CHsyw8teZWH0JLXoX/EaejFMerhvwI5iOuaCeSVDiRiFH8+HgW0a0/
JVbtEDhr9xuY68x6zn+D8LVW7vkx7aTcCsnwuIrVoO/M4Jiua1obE6sReuVh0fBataGlsZRDO8KB
Tsvkw4oiI4do05CoSFz2BpGL2mypbRfNBVTtzXgdzA57ciH9X0VffWHutDvytPhv3DRoO+T2mHRK
VDn4pWWlMbdN7MUI3pcP6GHkRJCi93xLnP0Kz37TKFkYQPfGRmeU9c68ms4HmDtsz12xvlZMu7iD
Qo7FNpyoyBoVPKZPj+/hieuVRx24EWHTMF6KUCXyKXwnkllFis7APTcKGd4SzB+qKu/aNWjk03Vc
tIKq2pg5kvO+WngFZ/jqrtJFBXWgKrGuFh9/+ew2BilXBzEnBYkNIov935GbAZIUI5KlX0e6YYP9
eK03OW4cYLEtfSqUkjgeIvu0U3uHKliVSPEvqRTMj//CNVOhtuoZBNOPEvrDDvEDNwh4mKgqFhS5
r+VqLl5D138iVI4ptHOjuLscmFnu+T5vBjaFm1fpxO7MAfr35Hz787JfOXDmLFIkp7WP1Ao+KpIT
jxblGglB0bdkn3Jx3u0jYF9YODHP8xaVcu/N8FkXoCl4yjiPC2lm6VknRspROnWIR4J2wYw3/7eF
c1AO0Fqte49RkqRhpG0v2U0CJLQLO7Q+X4LPVPFnPn5BSf+XC5zi/+LKD5Eko4MhxHT6A+feUH2r
Rb2JJb6zBw52x3srjkMO4C/R78n+mcWb3TS5q0H3VjAD4Qxk/8W708ILVQvCGXryFqQCCDtzu5/4
6mAtyMbeHiqfns6ZKiSm0DpMzrqniwD2H4vYw9dn6tadc3NQC4IkRXWck4qKvqxT7+B+g4KZ3Wy/
SsSIqmuAqUTTLuxWW8DaJ72CaLJXYVALpXAS90Q1dT+NXoho5bUhtMGSDo9WRlk38jzB0EMlxItx
s5rpcL0pruVpPBhPkOoQg6JGHDzmRLC0xe8a/C3lDjgLg4MVt9r/z1W8KKEl7qFIBc9HJVH8kz7j
zFC10mkjH7dtExukSWXoG91tX/AbbQv/RrRJltaL/D8TocQDc6wcuCzVq/NzZRmIq0K94pWAaQSL
PUGfISWwva7f6JW+3uoM6nSPb+do7wokuR4k8rozx9MDtkfYqWYSdwmC6rfLYnE+XTwSdgUUZqcD
uwUKZ3QuqoQph6lGh6lNkJcD0ppfARQAe71He3sbDyV/Ur1uN/O/EEr2+HKqKUtdnABDxRFE143e
UsmaakrlkkiSoIeH7ss9V98aDHVMqPAYl3qzJ8yDqbs485nuE7zx8LHh9Oly4agtrtHlHYzLTrBO
Lt6Y2Ygkbm3Y1zYm63U0djrfqH8CNVMyXfIHeJKv+5TVPuN0Q3srYh//9KBPotyb6r0q/aRJSZSR
D8vsxVYAWN9NUJq5d0ftRJrb6DX2k4cQEBvW9P0UjocsEnHLb0u8txFFpXVF1S4/94xxcSoqhzVI
hb8qZspZPyCfpGmSaOPceL8utnniynPCIB/ewxm49nQx9oIJ0KQfoTzdDpX8hTpBdkVTjgV0xK06
RhTHFx6Lqt0AJNR0VKqGnLf5aPlKsq0bEbn1I8JhbskcGeUcnBpr0qKnig0jfodWLKHyOBzQ3hh0
U8zpWvUG3uLRMvfe1wVqXIR685CfBmnp2EM0EE7b0mX9+cFctq4DIJFuX+BRW2EEprda5/VDXC8B
DpAsMiTwxEDmMpZg3Ak2VBP7FYZzyLQXnWz1kn9FPBMJk5ayHn4OVkB8mTrzoAYIojzy2/xKgQ+l
pQfNYz65bTXp3wulZJw5tiJI9Lp5L58z4Zwo4lk4SoH7BGJTZliwbdcA+y+ljP4btwgoYS7i3kn5
2gRhrLOvfAxp8krnsJ3wLIGI1CWKNrUTYdgvSecJM+UHpI7MdODGhWG31/guCctqOGFVxFOPVV8/
R3eLTxe3YXDwdk6SbfM1UextK7ktJY4DXRY5LK+rdII7uSknZRCiU5X4n3pC38zppnIEC80VLbVI
BHhmM//dEMNKTKW5G53TUKkIAxZJKnl2R9mStZqw0DulSKp5kkM8XcB/n1dhHLbJb2L62fpzGzcm
Qm1INUny+LPh5fGRXfrA0ykiUhBZ51RvCDreWWn6KcZgR0j0NdVOxSmYtDFNp6IVuoYYMjMxirSB
L2PHpxHPyW532PX32wd7lo2Wa+lmEGR7piReLf4hAvw5NAh9BLn7Ug1nti7picygs27fRjeJaQiM
uN+xWFJyL2SoEPUEcO+YjI7dW6pOl0t5CeYw5llJqvFqgCHlpwyurPY2KBLLfyUTqzIvU9V/vChJ
1h6MLL4owTr6pjA0C/tMiBIOt294NziWl4yOy+noMG4Z1gCP+OOdIcB8WaUsM/2G0jexdnqSXBf/
92P8jg28UaLf/l19DASlnROYknnrtOfQ2vHi1x6qe5XNjaMG8N32huaIuCWfNkJfCqEfJcyEEnil
K+UrXht1FZpvXqf7UbYSdHqCOZMRNnlC4X6kahH4/NFF5uFy0uWUba5CnLnUlsqIUH8RmpMsYjPo
N80pmDbD4d0WqI4EteX7JBEgU4t7ai4pq09QIaHJyxkePSnvkQCQT/FnYwN3cFTFKIzv2BvdXvWq
K7iCrWV5R01TGQNetBlvRqt6Axy/wtzGmSIXB7xQ1q7jKBRD38Fp8eoOPev2c7CpucdBY3OKxckl
3QiVx1TVcaaGZe7t2a0IARCsdx8VrVR74u9dJMwlA+95vadNt4fBikuWt9evm132FgYsgeOj7bao
YOq9fgrHgoGpOdCbiG30mEqaJJ/tzKtsP0vaAJsJRe2k8ZrKGdKrYwaOe76VzU0Ya9whLMqQn2lb
jVa3ZKz+mue8VMaXsHGwzMtXewHrpOEb8B785AqyG/trymJbxQZ378mkf1OszsD+dU7uHMcmH+J1
H2c2z8d3120kyBGhlQLQ5+5c2ezbAla4xbxVmNf9XN5aAIaW9zez+j8pQQ0dZxebtfSdbIu8vmUR
rwPYIpX7ID+NMYoFcReRq7Kz55GBRuUMc1aiIdiN2EuKUxYrm905Yloyz0sHZ0Db7wXHyS+FU2+G
fW+kSs2Wwyt5+jqG7a9yQkwL/ZgzaJJx7AoHzftsA3KNaJpTlqmSrfTkmHIVCv2FRDsYfCD9yZYS
sfm10621eaSKKbQHKrsGcOYj4sGpI+B5coD2nbM2aMGK1tEoIcht8vK/iSvgZCMwWD3t71bNAHrG
LQathSmvw5jeZuHOYC7MVL2sRVup7qH2VHEi7u67EPnq/snYkoZFFRQBSXSOenzHOArw36mlFbBw
2NX7ll77OmlSaP7Wdh2hjwMZSIZXFuBiFdEBcko5rAJXJZNSag01dkVOeGHj1UeGynGpVmLyldkv
BUM2m+ZpOe5uSAGSmQy+MYXvRyiK6zZoKCfAfNsqzK9t6XlAUezYhGGi7rS6lUMo4me/AmixT86k
E/9qncvjXdega7dETUJjyQNORLwPXCYOZtcJGuPvsrKbldi8SA01G9UFvlbQzJpKGwNzoW1JzVOd
m+Tvg9AoncQ5qNZV+4VwQSJc7q8GI3w3U/eMoh9SYxvRUe552QUoniqm51vqaNbgVesar5tbl46T
Dhk4ZNpqhVkVQDhlbhG4ahW9bxxxxc/n7GCZbEBmKh+yoz/shlZyQdyIPtiMqv768rT8yGvZn1mN
/2CkdMf49QbgxF8dfPDqo3I0vRmghFqWiABh8vMMFh7zj3pAv2kujaj0PDpaZM1aej5z11tnIaH0
6+t0rjR2x0jd4JZwhShXD2c+SIWG8+Xvc0cHb6Lns4nINofI6T89dEp1k0tTiZnProTBr+MzkXZZ
akFSFd7c39GF1YY/9P8oChmCmM1SXoinFfG29KvJYAC6wwg1E9dwiK0M8En+iX7pFHFoEZZwr2eW
Y46FQKLJga55MaMDVqbanhX5jkfrq7rqIygS+l8SZdjnAxlI7b8Ki7x7h0WlWhzsF3KkBOgDFd7v
klD3UhGxYEpdj3/7KPl3yc8mzBeUDu8Pc1XCTLd23im8kK6T5XuktNQcIjBNqm9+jEj6hW/oDuL/
Ej/NIh9zhrmic5t88ghdXK5goSxzCzBnRnNO7jaYynyigmBoj7QBxm0tlqyfAP4Kd8CAPyz0U8DQ
y53Hr23emk5CiEVQTKUN8y3qbw/2XQs5rmwKFWVmcBlEJ+nngvCF/w6dTIgX/CP+s54/qnhlO9HX
V2MW6zjHQpsUvH1aSMfeAl7CWLUEHPkLLYJUbk7r1i0ZcLHaK1NZwBTutk0KSUYXZTh+UvR/jlMD
SnK0K6PFDBM+sGsl6RduXf9SPILhlU3CSxiS+xfEHDrJIV05G6i3Ztmz2AwbxnZAV/SZlznJO4Ml
Bb3rQnpFq/Z77f/jQLW7VSaJyH7IBZ8PycAu0av8LkX12/CcKZb3WQZTw2QHf38cKVuH3nmvgof4
ZCj876C0x+5MXmKDZ34xShq8A90OPfGWXFgCwi8CJUgyYCtgYJvrYc7HCBxdGRC6UN7kYKdGwhp8
DunWIETbRX+GCTfp+AzTH6z5ZhbhxtiXKMOSqgAa2+ula/yVwguHyfm+cxKwYdc6HbJrcRhxxDQV
x2YJetnpjpIeDOz1SO3PKQkGhKu9WOgCNUIL7qsG/7QtwtBvVQ5cLJfKHgueKoDHqkPPsG13N5pE
OG0Lbc+Hqfza+NqhXSskwhpL+hpYlCeQC1nVKTncbjbGTMU61cnYFYUXDulXaBF5g+nXMAln5AzL
gEOhZhEtxgmE635A2tnpsC8Bj0ut3aKucU5R+l66pqJa8inXdDlOCAQuKptYtkCMCMOLh3dmPUTI
VsQVT2Vq2FLPoBQTe7JF4xuLI9tpDiyiiBeuPsFznbdPLsuYwrI0SAM1mdhLXr5aIVrGORC8CmhS
t7J0m8uhQZxpFF/0mRssVr3y2C73CeHaLRI6y6xganwotc3+i5sU0428pJ3NuYCbrnhJZPlV2I/V
TUgdEJljZBKQGYlnQKK3BsSyNEkpssklB03usPMN7R9NQAksEzL+d4kxyGMKJpoEKpM4R1+6Yo8+
JWe2sUG4UFZmpE4Nc5lJIMiyLSTIsQg4RBAGvuGGW7nZEDL+3Iv5iTwodFN+Qz3/sXuHYoWO5bG1
MGfxDqGvq+ulnNi1Wt+NxFy1s+0y+YBDnkvYVLA5HFDY6kx/N9JohrsvM9ldMI3JnmIqWyQMHUvW
snREi2iZ7lU/EcPQQhvxERrB1CDE88UN2yk8IK1LSm8d2flU/vXSmFpEBycWYAImGS97ZN66boef
v3ysKIl6slyC4PgWuJvbW7x55oXRUOSRIQgeKeetwdoHOSwvmLrTLrhYtTujyruCHzCupizUlhNM
ByFRWox9XEps6aa9axsmv7aV1vEddwm0a5mnjfaIH2PzOJYYLt1Bd0CBb+ueHZvInG92H2iM4jv6
UNCmXTj5dDz67FNrC9RhT+G9Q75b/01F89Ip52oxv8OYTbHtYyZDULyAkg2IasROVy4YELjWSIF9
fjGg0U/x1SUnNBrxYv9N12zsCNSqyJITw5wSKPhgzXu63K/jHbXUyBuTQUyLABi/Z4OToar2RaUW
8DJtIAks/7BeV6b3nUE75+Pij7ILzxxy+0yuDvl8DaSrWtSC2OmPXa7YBoqtHnDkF9akqmoXlkHA
V6PUEUM8H4DkZuzAWRDWIWBf009tQfr6DDCdJqZuDbdDEiL/ddBqATTajcfThvcY6s1eRIe6Zwo=
`pragma protect end_protected
