`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
I0n7NAh7lPD9ghjhTWY7q5FVi1iLeBFtNrwfbxJCCTGbv7hyrzRl82B5+WKGS0KB8dT7KOh5qgE2
LpTWFkOceg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fUGxIqWLpkp7p+hgpMfaT86uYBfXa6tnZz/bjWOgnj91tJIjZ4HMCD4MAtgfmK0x2Xpe5Wb7NLPO
s87MSCVVCBiOA/h3SGBbCl6+SJr8kvCbH5F9/bvYCmN4uXqxsxbhKq22KWEHZToxndnWcctbnRQn
35ocXUo0D1o26tLxWwU=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MiaF3K4Km1PZq1kKcMCaubE/GNIkpr17yqdcPEkVH/mWCIEANuarAwQyZdqvJorYhunwizVbbQFD
FjZP2gz8WOcBuMRfJrrCVkBMcbBKnquInJyzCj/0qVbPulJ1P30gFehdTHRWAp7lWhez5WUllMuk
kUnBmgLdkb/EuE+DmBm7tyUqExPjQbjgUljP1Ut6Yd6swb7QD1OEJ1wk0BEopAMOueco4FaEcRml
u+POHgZQALby1FcEK+8BR+tXtedWu0DLDAjLEiI2c8Kd4Us6zn29oaATqNYzanhrdYgTSOwM+PE3
Z+oqOVYKom9pea7iP67dNwTYsbLLWunrz5jsOg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
spgx6sVCkLoyQGrTVoM0LLggqZcOWIYUTQpk1U2Q7QSZUxoZSlAesqGt8a7ujG01ww9BGpt7ArAD
LVZh88WY1tAVX82jnKzh7QuPNMfNI4WwKVkJI3CiQzEusVBtQ4M1fPBKItUzEvyA0+QUtTXS5Rp5
G+LLF0CqHqlsxQBWxABQ0rpRc1NNrs8ktfDtO5o8pEDRUcG8mrdH6sSlqnk0PDzsti92TfgChXf9
+P/D7KzGFstMLoTdavEG+fHKAnHbeX/Yf4LGHm9pfqyNg2pTGnapfa8vm5o9UMVCzocco9WSvCsj
doa+2gFH2v1jFtXZgOh1Pfinpf6mNIVEvrTpmg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
l5uAZd91bKvtCPTGfKStVfJ/YcQwPEc1QJSpTy2G1IZaFGkZ2VuNDR6Wcj1roY27HhOWV8Yd1whL
/f9j1AntqRTxMpfOkX8XdZZOONq5w7+Mdp6O7eRbBunGuCfnuTq2ysecwCzdBvAWC3VI2NAs8lrX
3mNW74wwKWzhpShZv/1T1bC+8slNmlm8YHeC/5xvRaIPvXewkTQ5WWQEVQ/WSutnuy/3/ZQRbUSi
PSsS/KRuDp034MGeSvQcxDceYeyXqZjJFUua1j6rww+/8pglaSklFowRq29p24zU+8wjQjvRveC1
HkDsqQScm4Qv3f0xsoo/slaciZypQ+rDZ6TQXA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
c+DB3pUEAuBFXd1H3t+yms0J2EMKNwI3jBYkWMq+YxHY4XgO4QSU1vC1CpvU6oHyQk/h6yOgD5N+
V6eZb2aAuMa1b1aYdeeo5zHszJZWHWuSqw+qjw8iD2wuJ9lZ98W28ZVvHcbcJM2MZ89WJ2aKjKba
+WosNIUVJ1mNKhv7OVs=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WCYIyMJb9GXyx3NLwNdDRIsLlZMjmFag8BCvf+pcuxC4FtORBfd/r3l1IkUQR231iCqLPDCl5AMF
aJcZKwNHm0YYti1t4+5bKHmwQWRPa3J2D+yCVjH1cV1BuJazU/xZqaemQPB0dIgFfOP4ZkbttE5I
Tg5YEN4YAPMZAhZN6hyfTuWiU8749sHYa6d2Ox1iHm3B5GyU6HOXKXZWg+UgbtVT7rR5IQecGZHG
sbZ5DpjlPLob0w+ctwr/o8Kmn/Jo1zFIpCXnBIaVUVnyvAOGE63/K/W66tmOkSYxwF6GIUoZ6kVR
sPw4+MrbxZn/xPQh/DOGe2geS1PV/uZrzRQSSA==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
wISAlnbnTQHiY1JyL4+OR/F6r17CVXaNVzt1ojURbmsRII6P0rjnXmQi0pHB9nDaMakKiQIS/6jl
a/IM7qMNhC4rxshGk8FkR84FiTb5kaNXnxVRd+DjcQr6p2kyBXYea4u7oUQ5Wsa4AynUfNe6W+bP
Xe0mC8Dfpli5JCAIv6GTufCytdIF5p61TKUs8eP8pWlSq0U1tzrriS28H4Cu6W69UK8KQcKCRLr9
8Tk/ggkLrbs+bSuHBdv9hGyyNJi0WZZk8pk/8HpYFFoTNQkcfL8kSDRMNJvvQRmkc6UVwH3zeE3f
ki/RBQIhr7A7610ZCWRBAVGj2EHh7N4rKw4fvg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135968)
`pragma protect data_block
EfreCivSIJjH8rlCp+zLAPX5molEG565xFicuIc9iMRik86yt/s44rc81so/RRm6h/FZDb4urn4m
YdT5jMEPhIU5Td7TXHIp6CR4hpH8sZKUdBfOK3iefajF1bhwqYMFtRyx9M4Z2ukkfj3+A2oobEyU
Ju4HG5C0cNeZWP3evg625hngGOaQhGq4rTucsBOgr3FSOPlTsdIAFS/9L/O7/PwDSvZBg01n43Ex
m8hTtB24OKKUd/1t+Vxpabk62GYqXuw5hWVF8r8FSDDZDC9NJ3pQrkCSyU6syqGKn8sd4mCAtcyG
P5un9IHFXRGx8v0JwEoOCUVxToPFV3GAWidMZXXpPN680ovbD6fuJiYE7FJkn435rx9u/GXMLN3L
wPgYjxxu6JymJLPE49yUppTn8CfUUqCWviPMy0e19amgcSJWF3o/trEGDZ+sqhJwOJ8UZFIWv4Yi
ZtwFgUEZ5GSoRUrqpV2z2iAH8lvoxbTDXb82U0puoHvpT3C/eTjzwIhJGGbGzZmJWYu2m1oqPT53
5BOm4F+6NP/UQ3O3Fm9ce/kKDpw+tqKvFOmRwHleBhHheN4GN+6YXS/7Ub4hfg8mHvSYJxA1HRcb
XQ0++L7smCnYrqys5dC9qQAx41jksYaN6EXvvD+4yXxDDje4JnQwUYjYc5m1pbplGiY8Ep0f5IUv
2gRr0iOJj3CCTcOo3bEttBOXtba4hGkEHf+eljuE7dXVC39fb/YroEEl375k0bPutJ5Ty7Riv7Kk
w6wZJVU7QBUdxRJ4wn4QUmu1qBcV+ploqie8Ny9pGW6irL2T1aYEuXE8pDFslT+/RrOihhqdilz9
zJBgeIemJktzPo/NM6dsJn/96h9S7UPhwqEc1uuKK8kWsGPHB9Bkdz8ZU9el5X7OHug4JtbmdMzn
bEXPaC6ZkL4fWv1zt3w2AD7Y7Rhk6KlhKpLKUrnBuCMwMPluPbLyNGrXZDVh3ESOtr77LVz+nYgE
IA5fUAagDbijgM59ShlXctImbfJE1+3zEJc5ndEp5wJgGPrW0geLm0pUAQmkbupvAZAO5kHs2Qk5
pd5gH29ybSxefGbcAN5tKAPrBwuBAguWvl1BDt4zFoNdt82kfyxB77oxQTs/6IoA8I8fPRFg1vXX
tMdWm+2r1D75BqfkpY/5twU9Utj6lX6CXJKG9/VZcXEiE9O9J6sf6euaC9f2+fH2Od/zUJdEyJ+a
0JTiTe5YEzXJntPeeZ+SRdN0LPExjq8RgYdPQs/pOLkpIRjqtfzWWivZ1kzavYacdR+lIU60I9Yj
PgqEjGXNZBj6U3p6YeGG77Syc/jZhz0aNrQiC87JisMqK5b/6XflXu67NSbvJDpE3M4tsARshiPg
NpkbjnzVp7hb2ImvNwgV3ttK49ywd39iBNuRE6J230kvCgeGuxXMPH/oz691o1S3gli6CZS7GVc5
ZlR5nthpNAxtOxFyan7KlmNvNbG9uad5kmEPr6Pc862klRCWDJVBbOTMu4qEXCsbYnyzoO+vegc2
jAh+fBSwVBYwMZrC4w2WZPs+EGHWpQ01OghEDbW3rXoX9U0Svgr28EC8cJQWoWcJd1Pb67fG3SfP
66ZSxJqISHo6LVL1HdyKaKHvufDXkbcrKPFdh5msZw6AZFljGoTjBkqPpg6e0py/SNBn0/Bn0elU
TA3efHlSmFjtmPlLOI5OlGL8wKV+u38E1Kcp9p0IXsitGMbp1xqA35itF16qiwYpU63z0zzgPusR
eoYouU5Wf0m4h5JqrPeJ704E3Iq48BP7KELJDXZ5TrHeKEG46nVjk57e6/vvkX61BZoVaD0Giz/+
XXNPU5oIlBvtdIDt+TOFKPJD2crGrRMbEBdD5TwVcceQNRx4ygznnJKUmSwqeltc5gQ/FScUU8J0
zNb/yV5x7iPrfh8EYqdzTogSCW58y7XoYLGRCY9zcFc3L4xyWKzslbMFLeyNTBRD9eH8jjvSbmSD
ibvzmIFfhDx99mM9Cvsyo1qbzZ4iRFHccrA9BbVDtqvVZPft5j7o5ccZhBQjo5bc5F4pogq9kWvU
S6fxrEwjgU1IsChnw4MOzrT0j4n4Q0eWBHzXGOq3vPQnGSr7uqqY2uHentCl4PcvVKcAOgx272BI
N0S7qmsErNxRBJhR2pfpEbwjEPcQpGab+alXxI2Y81ovesGL97nbRcqS830IHzzLC/3ytcY4rw5K
LVKmIjqZ0mqYcYtAfVCO0gEo/P+EUH0nwejvHLnVNRLHcWhQN2e2MW0yTYs+3cR1KcuieWKmKp3q
HYbcxS6hM+z2dXWWfrUHGN5x4uGKfxzmiHF0NnKDA0DearlTYPsUekigTG8+g+yZQEiv+YKIqNRc
SVKNVG4YiWjfNVZo1/HozOzfaNhp3LUmaZk720SoRR8LiarHGpIC6KeRoQv5mS85m7gm4USbOgR2
ZEKrHlH5nOuDykvEM8e+gB2vHxMq+QRbqWjIpyY6kIobBS7uIpeMAEWMwq9NVTD9SFM5/9O8qOfg
KRKlyzXQmLEEbtHDd/Kb9KC8EfcjK+35bwLaSqmVbGRVMmJJtb5lttCA41zNq4sUOKEBAuG3B5uu
6DK7AnjefX8B1axh7QQl8odlr+mIBpXEWWmULRPoFeP74pG16t+JtLYqSVFwcysCZtKZLNTTti42
FxbR6tvM+8Gxljdv2VgzoX2+S9Z4H2/xiys9xibJvMWwID0+CdX3MYL6KATo55JQqTRM1Qf6+edB
DX+yjy3L1mijwoqGNlE8zojCCN1mkkVQ+Ei7rxWthhRFEoUYWrZj5nVvQiZNtnToh+j3qC27n7if
AiR4lDWQzBvkvIcJ1zXyhclm1zjAsPq+kAfwfvsYp4+qVWH2r8QTX0ZrKeq2wdO5VqhEyiH4b7bN
WciTpsicBw4njO0wjIdhc51Mv/DGD8To1IYzHjnis9BD+Pai8v0nfjA/NGhhKPSqq11HFVwGxvJ3
xT+cNz0yCQciDlT9Rt+nsF7PQW81CdDycjJnSQoFVuoAdN0Ar1qz68+YarFMjQb4hPQIBMdEA43N
Xbxxv9QfOzPV14wryzRv48yzIHKNQUFt9ZKsD3WSUYKFpCnDAnqaj9YxIZefs5NqXD0EgnMld19Y
wuyEDI26kU7+pdh6QO6PSO0Nw3qCoO0mWoKtxMwhIyiK/WNdowjHIWrxZJ93LiLVg7SX1+ngmuvO
ViLL21Fi0gDs2of9zyCU2+Ff/czUnpnWEsbi7emhXaMIw4T+whBgIZVVXgN5I20dPLpw+2MS4hyM
xkv/9vwxQE2j/RNIem3KY0y+MpmCJxWfM18E7DdEXGpNdUkZz8pwKneORWYkeyBSPByR4fu0I2gE
4pH61wIt5S2I1dt4SULChgoWf4j+zlJuv8tjBmVDps+WPSV30xVu2/iaOumNjRPMkDJFpHrwRRQe
c5zgYBdXCoKQOhG81fqYqDXpEotWmA+IVvLY86TkqU3c4wIXVNRvbYXm/YefjtFWxt6/szv+sFBn
mQrPzHar9ApY15jCO1iNwUi5xxrFpi3E0eTwVl4AN6DXwsJYR9p0apAVuTe9+ixX65R/8QXHQh+Z
j3uKtKW+Pt8B7xdUk5V4Nc0D8ijciLKDsrsebKpyR4bM5qWM2e33VqGlNAaZr66f0+1b7hUvJd9o
1a4vM/ZiGcBzjNMBgcpotldxuuIBnGW48mEqse4UKmCV6TbZXBiBQ3cHPE/J7RcEi5NAldoOjrd/
TugZjgBEY3Uyah2ug7vt5AWV/+LyR2Nh9eoNphFRO3Gg6uNqXe2GVv729Q67IbR1sdZ4pZ0X50ly
+8QBLb5GgwD2b7XeIQDHn/VbStt67Z6+mggHSTEVB/IgdmcCWZDl5w95+2yh3Bs/X77P7FH0ZTZX
xcHeWJXVitinzg6n3MKL2aPaEH7GXUQ6bbBw3JeE9e4RBhteXEMOiDiQVhB5PwNFBQ0sLwL+aByS
LpW4WMoDBWR0+9vA41/MSY8Uc0IAR3JzbZ6NUhUZ/l5nV2IaOogXAgXxzyoYQSepRxxz6cff29gL
fc9Tl8mJzxH0xglsSgSFf0eakJ3V0taTMwMOgPS5PjcLFM6dw1N18/IAazMO4ziDO2mPGRz7DVF7
Q+OQz3agln1IOEtslInauvWb0e6XdLN9BaztzJU6JRNnQBBk1Y4cJqroeP5ez+rKHJnxef7zbyY1
SSNJoAbpaIbCmNbjZBBnSC7RU+bA9dt+4Sao84CcccICNabJ6r2mOBZZCSgANF8XN4aCH4ypuxIu
Racz92n99QfMIwNN2LxXnKFvcAJwEOnBi66aH90eCdI0H7TuPwjAry34BpULtSEhlooeXr8whYZj
Ycl3TFUjCWyQSbjvEbIFzeDaDAsEk+wokrBMNEl8voGc5ONocrGlBQr0TaacH4fC5DmOXzDroq5S
EksC2smsK6I/kGwq9jU8WiLAS17j2/xpJRwP95M0QNLSC+gcUhRaJxuV5EBlLfnRA1dzaR7Blfro
OjAlxXP8LnmoKYvWUSkPm15iKI4zGI/KUO/xKgkAKDDYFGi9Jq4xi/hRtPmS1oixnIaumlHgcLQs
miAyGdBJN7ItaDlqyZWpqqO1WX32tZxyl7tPOUrY31Z+4+obClMlbMTcYr9WoIXtroFeCUx4FXT0
rrKa6xPJhSCuY509NyLI5040w0Grr5JpVmQyaFwZ910fG6FM3JiUiH3DX9vjU+9LU0DdBzmykDb6
8BZ5/ORyoAxOOQGsnyNWiZdOpgI6bSflXOKq8KElVtOYIP5XubruXCcKxlLCQhSn8AsIN4yhhdff
8UqQuxeE6IygZxsj7mLI9dbnLXwmVGQ37Uq5NwmUjVNnvb1PAfl7bPT9rUSWhfoTu1L2VCOdHEHC
ryeRsqOVJ20Hs2DSzYkHlI4cqyr2LPl7jFYR6Fwk1tiFks1EuKhGjybHLq5Y16s2EFavYFvZETkC
KDyIq5r6t3oRniutvXOauKimHBeyDvNmnzBH9isv2NiO6IIyAhd6DZaJnIGbn3eVGiwLQQL/KAlW
/Xh9TOWgNrSFGAoaxxOivJaCmoMsG15noAO3qq36U3hYYdU8ye6OKtqN7Wl26hlu8LUMTMOqL/X8
QFkeAzBPChNCGwM1snGoNulFRxAxzDaKAAqR2voX6LhVfLyFIXml+fmZk+ctraQ8tmeojMzXec+D
XOrIpZWaEbCpVINdFsqKmIFCpzmkRlEqSRtmAeLPOTM7S4Bs81TBlW4SV68W3/8XEO8ANgSZyo7T
9ZWyJDpJ4vuRoK4Ax6G+WUuWKzYY4HG7wgmmYkbq7pJgpGsrWZRKjnyfOAF9qe3XtUGihyURJ6YN
37x8EIRh0QLQfjgrN4kh0b2isnHDgkoVDVYkvm1kQzvFc44mnaaER4sfPDLtyxGV2XAU7TI2TTyp
H/cTzEXbAX5TctStVfCSLOiRufV5LkFUZljoG6Lt/0D7ySUM2AcPcFZ8mKxgWgS5z9nW51wX8+Ht
pP8+aC8sYGmtIcLTenr+K82hMcu2BxaPkulxqpw1FEjXtt05Eu/yRAE4aFxG7M5ipIHKht/hXyJz
GZgUCqoClGTLHrq3qAd0oBhXijYQ9Q2WRdtA/IuIvqWJBzJpTfz+QUI2qemKq5vwmbih3CMRNRaF
kOXRyglHGBU8GZ+W2iQKZk5wDjkViYhc3jxaM2xAbRpEjqKuE/7JZSb8NLQO9NPqIBLch95gtkkc
hJPgEbK78tkwIsk/Z7XbVomzR61Z0ADro00agy8Ja2uDfzSTeZF+wU8kgwqGnlDz6bZY6UrEwoGX
OeyKNPF1DN2/Vl8s/eTiSrvVPkdUPWkaBEmv40ivuHjdqBKJqcJBKDnZRiEtDROB8ZvqD34In+3h
qPNRVWEkHIKEsNFPDdOZXCdBjUjHX4fzQa+CzINV6Kw654WZDFKcugbFIrnGoRWYtb4IJUgXlNM2
mumoazDBOO3xy8SNjAH69cJ1n55KOWHBpS1rGoXAV7nm5sSNoPPrpivWDUsLj1yphdM4FmMm2tjq
yLiruI7igbK02jjbMab0Z68BTX/w2Uw3DT6sI1TlTAu7+Bp5qVBXEGGdSZmG71q1UFjs9IbU2IyV
0+CPycL4alAW0dF5vfjD1Ti2CX+A+GCBKFzIlLOzC8RRQqiuSHs90qkuD/uTFX3lTkvleFGO90em
iuRmI6hCGZQgA8Dj96xp+pbEMzLHI5+3fOS1+xCVG70S/kdRxMys8ZP6Ks99qcWuIplNUlfTehAc
haA8LIzQyhvcV2HQHvhEdW9WRTQmvkUyZWrSZ1Y8jdw60WAuXXDlD1DkigI3NTAtLbQYYdl+H0tq
CDhP0fopQzuSCl0i8yce+SMZBLzZLoj8t/0DB9VaTS5ttfqrsq/VlPMVuzfo7VoRcM+IvXVWsMbt
ZeHjtXHe3yYahbpn87yQGAUu6okRBn79YzkSwIfWvreREf9FTfv8YHOUT228oIs5PP4hAb33Wynd
1yfsZkS24Ke7JnlefqypMtv/nqO8s/37QJzWf5KblklIP/JEM+FkPn+1+RmKQamP3N/Y0HSK0vr6
gTgsepn1Xk1+yE7dhzVd8kEhI5NrHtUVH7vLO4IMKCycQUOB3wVVztoqtVT90rC1uRwPErGifGXl
Xult5mbTXvAp1veJ4Yp0bBNwBnwb0GTW6riJGrdD6i06MgWM3eWoUl9TYD+n+lJjjZ0Nx89epe/F
xVzLRtp5YQzUgWlY6YtFwpXgP9KpGD4f7U9/vVRXwZV6GYRIGbGZYxKpazs6YFRCJzrfcWO1AsHt
+1n21qyMnG+4JsJRIMFwJu397GsPKQ4YQ/x3KdV/drj7WYx/PbsVsco7pPI4W54/K4UuzJFleqZg
p+z0UYU0yvQcISQN868oITOvvlpUkP4Jlj1NkojUlrYzFzmSzRlf98YJWzndItTlYhcR2aNCLHwB
+ijMlYLAcxCQtQT70GvFHVmQz5Cmkc17nkzG8645UREjLwCv0407yyc/CCYM075KMcT6sLQugK8D
j0O3zphVNncDCmli6bargVISQODMAbCWFyFvnMSm3yNJK3EmE8IbSL1WKEznOCfplNefuu+38EiC
yjTZ50Pz9qZyr0ekdYKW9D0zjHFs4jYh71d2W7hWnuSE/2f/5bIqaIIWKlzl+wjyHKdYRvundfca
gtPCjo8r79qlePqWdT8ZmkTwDX3fhhUZCPX3KwnAvQYjBE4Gm7cle/ACAbkfznRldAeM041BQ7ym
sYihwkaW6c47qxAlwhk4AUtsu/+zrvNZWxArYh9z/bivecdqPWs8c36gDyPghaF3GI4Pue1bcS43
qAw3xemvkOqdR+mUNd0GhFsuDKm+Cx9SCjxtIRRm5WOuv+ETTXgQNcbk9zGK9OxhwLuNgBqEw70b
TWs0upfa6nOl5NjCUJOzJEcPNvljWrtK77Q7+ITOzpkVO4bHY1CwIpsnrrkFfU7PSZ3pUrd3SizL
mh7nX11JdZi8cD4SllsReK9c0hWj5OuVDIltY0BQFxOdSOLokGvPvwvoUqpEKdISY6a6MJzHbYYP
9SSG+R/zQ9IWN/f303eXo0uapHpQ+YK3xc2yayKsV7CJEkGmat22bKme7OeB6FRO/ZWDBy9iiYZw
rnC43Jqw3bC4RqGY/uuY33T+Vcx5tXRMhJVvfWMQ/N0sG1Mzw9hSZKHBnoBNqk1CR5jUcOxNQXON
+zMZYDcMmZ0dudKw2OYhs/fUyHI+htaQbvkI5mxosO8t2zOJrF+SyiSiN0TtAjQRVfcXmGLU/VXt
OT1HBXcVViUIDYj0f6zoLnKXQivqDPRVKdeILdnHR6KYL5Dv4iPWBucWzUMxktAlMLPuGxzbXu9v
Vy6R5hUKw+Eq3Pe4OP7nqKRLY2wp9owPIpV0yjPAdYKCh7dSDgNWpj0meWG8cu6slgZjSzgx0/ej
7Of1vGQaROS/ysV2VBd2cImH6ntcoPO6TRjnpXjI3jXG5WgR/W0VD61Z4d5kD3qj2t8rHtoBvYFa
SX1gWc82leEgf/uH963Zo9m/5H9PLtyFBNnH6ZoLoq9EB9r9oClb6FDP8a/AqEJqc6x4BKsRGtz7
e30SGkVr33l965wox/uhB6lZrXEl3KfsDju/U/SwT99NA29LQh8avEFW3vPn6rX2deDmcFwCQUxe
nOH5SRykgoygUZnpLRActbH8e8PIharMnrTz9HwPUziGtp+R6blVOSfk8YKmCGp/3GNk/hsH1ds2
Wmz8gu6dLIFD9AUTA39CqTZqDNBdG/7iod/KGGpcntYIc7jG6vkRBGnYLgQkzwoA3xBgT0tcFoTC
PoHaJ02PVhB0It5Ua7wM6DdcfInwe22tBxi7Bu3ohRW8NmPjajzKOZhH2QVd8Z4RH+/iXUqSFHsA
8lUM0iIX6hDuXK0kZMaA9JsegjFjQufdjwg1rjNv/z4M8j5bGnqMglBWl2q2BL8dIMHKLqSrPxEt
7FBybBz9heU02SbbeSxnRgIgATce0zjYewWPTiEsmcjNw0vVHl59PcLHFmohpTWpIkYvcAeJAC3U
Wx4CrBypOTSKsS1nYYmd97Z8jcdmTY+HZdKHU/bz4TdJMYNLsXRdDkoPlm2UIcdXptYttucSqNxB
VBhTbZgb6jywP2OrA2ArChht58JBXLsb7t4q0YTzP9OkPLMcCPw2PnlV5IUV2/c5gIHsC62H8qBO
FpbRPz4cSQofGJ31PSfrJ9ZmdcytBQlIV5F2gcBP0JvtfKdH8pgLW4gC5lATMWkBBOBR9ZcRbq17
DP+qxYXGoCSdW68FnzOFWYYIMDlnInLJ1pR1rJi1XjBvO8qUfqx9Ivie/IFGNZ3eaMqmudhnN1vX
XnXJeznPLEigIRSsQcaqzo5bkC+HFUw52O6zvTi4MyXuHzyu887kHxANVul/7nTAnYTd5uwXJ385
geMkdUakOCJLDK6kgztvpM1KtoOaDHknBhW3TJy56oJnJ4xbL46Z55OeYUF8Qop3eZQbUxJuUyWe
zK2csRrfWc0BB2Sr64PM94TWCdXiyWffnUxHKHtiCvFYdSP0r43OrPbHFgxT/56iBjy7nB6LnKqZ
YWV+OhNJ6uteY9Zyeg9ttJVGoSxUyENBlzMXx0i2jWoZT6B+WlP14ACowbtI2Fg1mKrTolHsOfyu
HwTx1EVo4EvmtDpG6vTyhgWa9YEZ1WCmt2HHtONI1tlOnpdWRZTSu/CvWbJ5MwNl2Fy/OMiHC8jm
cbN0yM9GCMQbc4fk94eioOk2murVNIbZqAwkXH6GgoDbY/kL31On7XDjpnudq4jYW02v1eMTDUDn
7tl9nZevgz9OlM1mpCrvPGPkpjCP553q+ESsJu9A6o8jxeNnzXKTw10d0Z2XZqnOd+qpRskenIYb
xmPyonxQQjB09VMHOb/X8hDcHh4UzLH2pIGJgm5SCktUZCWyoWdAJW4Bu2fBkdd/0FbWkEwAeEsh
C9H84RhTE7vjJVdJbpOylETeGBGekdsanRhgUnzkItCRTH4zxks/pwdADcgRHLfyHXQ0pWVap19y
rKrLY7TNkbIoYE1B5l5QRUMsLAsK0ncgxTniZwn4bcIx7vwJJ0DcHyuuEmT8FH6Gn8BCb2I3/fSX
XeWbid61PD1gJri7xqTJMGc+nOOgwChx4UnG3dz57ugZEWJoRPR0ZiIr3n/rCU8JwW44p0cgXj68
wva0CgO7dQbaZ1bZ1uZSy7oFi5avBWIM+PVdpOIJAvzczYgdJWUGM1Us1rJUGNHuNkU5RgCdpCFM
88K8R9IsOeH/p+rlaBov9pDIiWkGQiagmISTGtbjmv3poPoL8hyC6YtrVDPJSF+rrSIAa2ncs4BR
FC3h11zRMHAHQM4GfSV/aany8uhK3Z8897itDoXFeiIA4Duxhevm0QatBDoKYF+I1XUpn07ep8Gq
GrnAj/wufDAmUOvRzB8UmPxNODBLHoNbNw8iHcrBjxlis/UFJ1rQUkwsRdLtaoq8GuQUNaYeBV4b
m3CO34LZutaHYy2bLsVT1MThO0DMF9tMIVHhGWLqs7sUb9rOtW4lTAY/lDsOjbgVT9MySio8TbdG
40gpY0XDyhZqRDgaTsz27Ajl/L6zxSv5CiHSa9gxJIDPWwq2D1vaClcfWH5VJnjV0uRRMwOEQkAo
Yf10GHujmTW/uTg6c3ZuaoKNBdYt7xaulPaRDokYZKVjuw2hHAz/9L4yBwSIEdAHG6YD6Y0fj7Eh
eOGWqcOQoRcSTcyhMISNcLPEqcJOKp3+p+mW7aZtEZE34oEo+nYuoxBEs9ocHVBL+fZp8InfHg6q
AvAGlbgw8D/Y8GscNIpeWvO97628MF42Cn0pUc7re+bSdl5E6yfp/KiTVEN4nN3e2M1/EgkMUpiJ
+xKID7vmLUe1INZ4rUfgqWkEHIvyiWdNLqUsfyGAf7vjCWXyp/CfGEkhYiH13lTe3uKg798cq2/+
ZjS9T7q4IVOoIZZoCH8nfvS/TslWKzImFVWOB/tXiulVUk3T/+tcOCW7ZSU0zPad1b447SuI+vcF
zEzuQOfsqteD0FsYbYqKJ1nNCarR4Mv9VJTyrOs/tSK1s/0+oE59v0m5yrCPQAyOa0GQVi8KfRnD
9JiLSbQo1WhUvfN79/GDhe7gmqdC5hayvO206k+qnc2PYvXa7sAG74sPWzKZFKwO3nhDBhFZ2akI
TtoCMIG/5wX7+7ZiJrtFt2R6f+nPKKIB1NcAiVqbc7Nkf0GKLCVUHY5ufWq60qa7sBM5ORMTxBLy
oyL6NS5vNkiREJpqTSFZXoDqZ7dbFRINR7P2wRjl9E6rvd18fdfok7E/h3Ysdm+SkXpmTkUp1XLS
qReGWbYocpHNDKV/lML97hTIVXF6PF+XlkH4ocEOMLimmbwAaNaDdHHxMr3Hjciah4Ceqpfy6AK9
FgIxcHnQuu6ajRVe101PL75kSBkDuJspN5+lMOi/KlRXi4I2r5q69Ib7lDkzgLbWt092L2RKHLC1
gEymZZYYJsjtllKgTFBlCdN/+gcwk2mXbfoBXamUR3ZHpO8YXWutDd0v/vXLQJHQP4BNGcGY7XOe
1Qjw8/2W4SYqcea7v5Qvtjxa5CwjZV2XhOUJbT4By2plzfM46Q6I1/Uwh3H6v61j2XtDoG8J+6vD
nOR5f0AD5NY4naYs+JKKJ/ES21SYV431Hvu93BGp5nwdV0Kgjx4yhIzjgQm3xASRby02bYrpg8YV
jGvuO0y7d9EgJQNOxNqThNAUA1hC10XgpRDeTPAq9DLs/O3pSe3nlYGptp5HYa+IVIPPkr+uiJQP
9k04t723Ki4nSLdD0h6y199fLmk7Egx2P0rHCKfmnIAbQfCHwFktxzMMRNtMkSzS3xKOUIjRCG70
wXLSutvJH+6Sb+JFhYzknsmDHmkbul8ttgh8Pztp8go6gRvGPrjJlT462lpds4M9HICzpz9td85K
pUXzlNrg5AK1IAY03D1ViKeVCcM+wqvoxywYiqzKzu9XsDYML+ViMK9A7wu3a+E465/Cj5N2nqn/
a3fEmfHPB3ow719jBByhjyn63f8axMbjaaROfnLj78Fap7APtKR2x1VOZu5BAea+INJsAforBHNx
mc7RqAU/8CUNrsABDG864Tv5fZgD5kXVnoNvLRBp5XCiPiJFcLl8oIzZVzO6YEq+CsWY7HwOqCBf
ROhmh/TRTKIV2lEkXyAkbub8lvDKRZbs6WGVvxzX2csypIn8htrYtxH3jw6GCpA8b0W3XfLODgKQ
IpKpD14CUhcschrMyG9/SfijHT5tBjIJMi+kG/LrXDAchoCd94V01baG+P6nY8/TQgjuDzr32/Za
6QMCfQ0nzD8Tzq8ZMy9rMYeXu69VXGFbljZKPk5Ia+fS2YkA8adssDIUO9FM/CY1AVYD9ScQ0K4q
q8LyCaNChl/3KKo7AsPaX1Ldz/+G2cvROeTzwpp75Is0Dwc1c9VvPVwDrqAW/Q/eJIEk9405TUG9
JzMduueK0L/ODZuAw2r9qMNdx3yCBxdJi+BbdclbDWO06keLZ0RzwHY0tCSPfCTzycgTC7BpmPMg
0bbq6oux7xq50gfLbqe5Kv7M1wwgVqacpockSGkVRZcobYlRb7204JKdIzH89wJfYsc/xNy2gnLW
pBAwrYQYqcgS/ybx4Y2d6+PearDIJ/88flE1LsXIlrBURNLQ3fBlh878fSa7yru0ygD4QR9+MJkb
SlW8LbYP4igyXOEJIoWPQ1ka878+N4wuDaD4iy0y0KaS3LiDsOn3CR32nyqgmjMnl2F+8IzLiCDv
qe+9OajrRrXpU/QbCrQZbRbypIv461rbcvP/2uaUepGiw05ZXBw1Iibe5QfzvQXMl743mHwtikDu
nEzBlEE6miHC9LmmxND8U1pd9xr8GWBG8HG5s44z/xIrwxXkhovmkqbzt9EfREnZR2eRXaSgAUcP
kBB+LW1+OcP3IZg7qKNrCdbx+ubAQMP9+7nZZ76NFLgI4X4v+lUOSOor6PKYWsK8hxONf2N8pGN/
k8oViE0uFx3cdvpbT4vmbFmOc0fSLJ3sGLrvhGLSPT9uwR5cOPFA+vLHxXbWAUSaN87Un7BNxQRv
ZDquv1RusmlZdOQ9CW1HFgxC855fiSqTLT4Qm43a9GzXVup/8U2NqVEMpzbc6OWE6x9PW4999Oak
0RlG1NpVdEXGYdZyGKO58HFl1ALO7CmihIfPMD+z0BXMH8Y26Mrhh6TMUYh8ZaO6FVYnlUXrxmDQ
B7yxWD1F8NLRajIkRGoO9romized1ttvKsKnkohvZrZjgE3FzMeOYFgz39yVOUpoc3SFTEveg1s1
asJhuzgo5lovQLhsO1CIddsHk8Xh7Z6iWwee8I1AnM/rX0aYERBvQt/GF03gwX+e8tblBB5JHKNq
9swH3AIathxq7zZsn9AsZqHi6234LlBmp65wCWUKI2ktMhGvSicDBNusTSnSTE7a/zK09+LEbLMU
9KFKTugZTN2JCF4EJsy09OLoK2ozqlBAY3I52OeKCPehE8aGCJS2NtX0CTd2XS6SQukSlDD13EDh
G0MTDxsbDyo/HYe+Xa1j821a4pIdu5fsk35MAFkLcnFdBz62ETlX6Ei8d8HVJPp0Vhg77a6juQqy
ngvZ3ETP4Vr9v08fHuF/S5JKGP2iUSOR2AasDZTHJCCHcByHnEQBikFF3MdbCYCzd66FE7NkFxq/
E/NMSn0GtNOkmY1/GrgOiEJheNKPdYsWALLqHnrHmuln3W6gASjRMGMM8CHsFX7NShSGVH5IawGg
bCp4KlkBzCPTKGMSaZTdSIZaz61mBH8iK7I/A3uzwEG5seZbEgMFJs0rT4n26QB4riryQjT+7+RX
i+Vg340wnaM6nrBzQV5jK09Hp0FEdbYH0pvbP62yO2g0iIo/GwYGTuYkhuz8a/67f9tTBcnzfAZ9
/YzqITwTQGFerezSxA0lnPbexXAkr5GceFyqh3OL8UZdAuxP2vIO5V+Tk7yMfmgdqUteUH2h6fti
1ARyIvGR7uf5rM2/tLRCqqyXHKI6UUOwpX5oMu/VZtCxiZ0EAa7zmF5fq0PISLRxQ70++1QXNIoR
qEe/7ZmPnCg4Y/3r2PKBz6DpgF2LHtepvAdQIyC5CkoXO7q8O/XJydxjxYoFEgDKk7P3CKJvv+Rf
X7zVelJ2F/g9XXYAsiKP3+leyhjEPaNEnIlNECWa4bs3nL26aFk0VyVbUYLp/lgxaNXiiECNnrTC
nzA35v614NONmICuqohGpJRK9bzbgVE91MTMsy44XX9jtDq8uiotaL4BlV8NkrnxTvuw4K3yCp8l
hJxAfjUFve+TZLaZpsksDSDg5ln/LEJ38Gx+6W3xV5xcNj3BtZTpCBwmQ6X/flLhCdlop90vJd9a
BBFYkOYf0NQXM3PpExVk9lgT6rEAYs4FU7Wv8TEAnn7Ul9gzwfhIuceACh1ZAZO/0tn/5v+2tqck
yh4OOIX2+TMD6vWJYC3P+gF0bIkDinJE4HVgpvYZ4RH1p7El9KYiRNHeb804anR1fwN4Lis2PsAC
2+NrqcjIcab4VVRrnmqIxqKOhq4e7hEl629WivzrEBW8sbnyicR+bNyIAGuBJV6iDXoFkc491EYe
iY8SEZeyzP2+A68C+LRCsTvi0Q7yyMLRjdQNTqXfvfK2pva4NwZbBLmI7ShUifhlI14vs4g3Rdx2
oRO30xCTqRY80vT/Jb8dCBoYooDLEyKkH05O1IFzF7Yy5kHlrzwa7gCHipisXbPidwblvZAOejI/
slZhMjEbQxVwoXabKARDjbObmyFTnzo6RloKTLvp57lFr+kx5rACFBOMTg+ZaER55omvjcF6qrr/
d2UoF9rSyUsiNvfMX/32gVyoVkjehgsOMxaHTaoRfFpgIeIeW9KjMEVK6QWjKNeAmuqy9NspEa/+
ohUYIS31QpwU+KgPg/OgAOw1H4OG5X7uee7hpi+X6qrCMP8aJ3v9kE97A9adq0N4x61mZI8NvpB7
b54EEu/Ovfr6hEl7ft5sOdrR4EMrj/lqSMYVvDFBtgtZVk8oifeHL+ERQF6ey1wtSzdn2y99Z2e8
M4bdNgoSUDEtoo0JAdDjjV1vYWuDPMTRhaaf+bb+L2VQDydMrFL6DyzcDVbjJIG0yqrE4pWvlEeA
MJWeKWNY0LsZHBTpaHuoTEZxe/2CQxbj9F597HWAA8UZ0XWrvHmnXEeTuv+fD6M8qnIwFF/Yn4/N
TCTGKl/qEBNpdnQIcbiSPXEwXvHvFbdGnqUCx5FzkvJWxLqtJxsMWD2oIDp9FcoP+5ouQXz/loph
HGEftWUdkxGVz80E4E3Mrj5a0Ix82edvQXdUEWiQGyzDpoZvyqbRaqL4GNyPtZvNZJuVGXQJfphC
XFO1vTIWREzjGCnNiabkwY9cNYPeKtSJa9ShMLx5AY9yi6J9jdaw4pcTYCeeQSvAdDu4IvPn+gw4
quhJeuTRslSdQLFJCQW2gYTuGt9qo0C0MvzzCZWCUFlJWkJFZ36/BzQZDWqt0sGkSlQ8xoCdyQMd
d08LgJaQAy17qHonu8f2v1vXgh4wunoke8ATXzW6J9uoBbtGf9TVNEwcZBfqaVzhnNlUM9AmTAGZ
Wukzs4PlQEVudx7se1pSlZC5hFfu5s/P/+bSQevQ+axi4uPPovYZGd+7Vcq2j+tq2KqNUT3ft3Sk
yd+FnAv6ZCdEkrijzYhj2HOcpA6Lipkrxlea5GMKmgrQl/0cJLpex/8fMIW+YZPIntgky7706q/k
0uGH5VMuqegdXqIcZEKTjteXIrYitqqV6gFNw7QjWNMdKtu03pTqmRaHungK+TPJlKME2iU2brD/
5abkBVNjc7RF64Yag4YHsMvPhA0MyDQYV+akWSmVJWVEZ3ZY607N7SR/BDB7V0B4xpPWsYVakpKP
4qZLsWH/pw3vFC0AAyOrsWn6qEo7F/rvKIO/I4ZctX8N0owQWcXEdVI0Aa7xiYFSJXmmFDffJ1ik
4HhOkXw9gB5KJZyb3c6jEO80sW/KHnNhGjGIlGKDGDYh0nZCgs7NazPy9nrzxTw6dresugvGnSU4
g8eXp71beXfaTtqB7Y7aqGBB1eI7lK+RsmRTgWPvcA0JsFG7yskbNhGH4AfZetstREt7aDHRQCWK
g9VJBbZVmvBWl7kgJa+/fXnOgn5cp+TGICQ/OQ9xxVfSdiGKT8cxapIHrHdiVrMET9CMjMUpACC5
EtNc44BFyEcL04XJvMp9E71fUaAtoGqR0HYj0cL5+kM9xBGynq6Bxyy4KxuEUrdI5WS21r+oTjfr
OVEhvq8lOD1qp4p865G903RsgZ3CLoKeHYTblLtvuaTsc758rUHtS53A43upLSlzDKJ4tuaheA4R
7ixYpfP6/3wcYRrOdpE9OYV2vc1eoRUzaq6TOiWq9koV81p26IdLk3FqcNE8bup4JQY7/PmVefp3
crUPXFhO+ebgQ+XAalLTFaVk/6bCbKanYST0n/OoOrrVAshOkZL4+Yu/1oDj0qKPIH9k4QP9vlRU
7OtE33rV9w65/r+en+ZwOEPEX2t/mmR6PYZ3o6Uzu9ZelYzODRX64h5+L8c4ymO1Y60tVowipTAe
T3Rc2L+qSZESySaGx5BKkILer6U9FLBUhnjniqe7LF2ghpRASjACB1CkAOdlkHrY8cAVeaZzLf76
+2mEHEh8F7n48CHOLSW8eXBqSQMuZxT6JZS9DHJtjZ/6f+R3O3PD9UEWR8PeFhaU4PKg5BeX1fqC
B4JZBRXe2BBOtns901fPGEJhKDMizxRVtxlBc0wVWeCZdxSFx2S+lRLErki6pJUSx6ArtIlZOwuV
YbDP8nQ1DfyH7M2tEHRHVwhOwnpBcKDt/BYxXvs/c3k9ldK+HHavpkt6aPWbmsBpn94DFsRxLgNZ
CYtfFcvuyhpKxjMLG2D9nKPFuuq72GsI12f25AXoftn14vxkvk+IwCFe0/wtXGXdo+uw2IltD7j1
+dpQi1ITSW+ohTLuv3n5TSesdLbOPzbY5mJBPZyIBOboINcu1MmsY324quSy55QDdmzaIviuvoth
DfeujsGeekpkI8OniFPH9jVwt5eKTuszb2V+VxcsVW6tc0zx3yJ266gr1+FfpnHf2e4r7YBS4H7t
FoFOQcwIVQ+SxXFBKx6eox93Ld3ak75LB3SQtUYWNXk51zjNuuVow6o7HObib7NHi3xiU8VmgBeS
znkKZk2jW03Dg29rog4M3G5Qa6K8kfDKKkZYkqOnnXkTVLa3N9PCrPL8J6e3KWI3via4lWwX6cwR
GhOAyACJgibBLGfyAZKUJ4OA7s04WZxSkG7ay44qVe3pfcc4aJ0TZLfeI3t30aKjh4LeZEuFpw68
nZZ0YFfzIjRkLP9SGFasjzwrUgOpLrNIbjn9VAydlzQTVdNXf3GPzKwsZQtljCn3+WVQWAYrQrM1
GJCTc3l0XI+yrFEuW4eLvWEaosN6QjTqMyBB6tUpmGZRETIefG8cyAg7Ny3S3mjC/FH39pKgY8XC
X7OdeHCkcFf39Q18SnZYWJXD4Wza6K+opQrRf9ZhzPIcM3paTfKyVh5qjdYtLS9cv1g5ygEj630E
yqk7i1+fbmIdfafTANnO0jwWdKBTgwLJCwlcBdUB1XhU0jz1+cCMdMEMNHAfHk96tmtAqi3pd0ZG
xrnWABpANvon5jTAzKnWvFaWDcHKVZ+XtxFh6c0Byb45Yy0bxD2695WSN4IaW4KeT5pW7gfnd8yH
J83OVznAX6XTu6qLpctnFGWL6ORQZ3wzAaqOXGulT+NdLjMvFLO7NBXI0ZvtXHDYcnBiLYyw0JoX
H0NjbVajrPHBt980ZQNH+0IMhzQD+SDOilb3w7u9RjFgRgl/SPbzme9+1B6bLHdapNAxO4P7bjnz
2PpsElHpJP+4ucBYS6y9fDopD+9VYW+bArZesasCscW2+awzHJ8yP/70D+ri1HpU0NIpxx+tcNh7
Qz840118O7TifhCZSqkbKalgC9TMRP7HuqBBAmZA+hRBA9KvvuJh6tnsP9V5VtcXmePG+uW4t3R2
l4oaMlEZpXm9jXVgL3Z1UQz0k3Qg7PdwCJfJu/538j4/xL7d0pJeBevfbsfh+PkHyoHS0QTP2YTS
kJId1UYkNaXDdiMMl6zmHWjDu8A/lRhV8XjTVOlAtJKF0/xuUDcJei597t/P9yFHwdb72yxo2m2w
b3nDQhSQcWi3ZIEKikwx0f8K52/qXmsSXccUPO6hYulydSs3AKo83Z6e0PyFXfjz9pXl8bMps21w
MTj8GViFmlWJwmfqYAVeqRoP2/s3AWS3porhntGh8BWrf7aQjgZiT+CL05QxXdC3KwDUm68ybm32
x91ymryir3haaWcoJqJbnIzJomwDTPrdbj5nNJgc4p1yGeT5ssEvYSyyG8Zv+vY8d7XU19z1u3in
bz0C6BPeRWxWFaDeU6wynb9Tr0NEbuAhK8a0LClowpBrjDFEIqvZnBIwGR5Puhg6eNyL47u2ziw/
nORF1tQ+8zCXekJp9PTj247p4AVaOTKdkWJtbcTG+qADxKomK6deBnumuUCcB+AisWhLVJpv/lNF
EVAuQIdvXdkeuyO33l9hwT6UOkQb11cWcczH2L5Fy5kEWqaRwCYe9g+Q6MfLxUiKX8FvmIH8PWTV
ovNamSNrfLW6u8u/HVKtEWDdAC3Aby2qq9pDTMsD1UekrLBNmoPbFhZFFmBfm/KfgjRRMDjwxaMK
i0SHwbFjP7+CCT1E0/PAxn24DUauludt7TSJIvmFxLb6PKnRVNanfnLuuclWsGfjsLB1s9K9xIuU
X/yOzu3v3E3X1hlfNwd6SKQ65eaerZGCK8nzfHkSJbm7taqwPpOJmM18i3Rnh7TSktx8XAvEkHDR
h5vVTgCXmU/ruGIsMBOIWHKWvNJZVGuto+YjoC/aOeSWoDQgdc8mQBMGK/FwlucrBLdyWITlCLce
gYD7vlVOb+NPa8/wSjeCsnyvhAM5Dv1We0B0pPpruzGHqmGX87xYEN06hyUzUxlvwtPQAusLk+tG
nUF7/iEnn0k9stGZTUUkUCuzPkGeOrR7QvpIHFoOWck17wfqhgZg5LM+lH68FwpUFe+Pmr5wDoZk
8itfStXQwG47q116+Ndwo/Qlj61kzNrfvK4pRarXDA61OvrSmHcAPA1RgOy5loEmUfxvWMFJNlzP
uCT7kU5DDDWZPAFKV0x0y69aSK8nu7oEfJxXnkFKO2qI4ZDKQ6QCqkuWdIyxsSSpT3uxANUPTMry
qFan7qJAOReM50mEvQ72s2zkFFPU24l9XH2AdzTY81sKsEyUmryZt7tOX3iVao+H7kOT29K2P5jJ
q7BjPVaGPDQjrSJ/oLflH9EGdQ9HNiV5v6+1TAxeULn8w4S58XEPIq1KqQkBm7QTHHltFNKt3HkB
Gc2CnMMSqUSDfuJZQUmQJEDXNTy/MQW2GvJzuCEv35eiP+eu+j9atevFd9JORn4Kyc8ds2jpLJmO
zRzYZtlm80PeEKSoZrMTIrq6ZY+SNmFj3kjek4VV2va35MrKTh9OmDmTd7GhCDC5MS3QXcF7yG2o
4m0Y40tpqldnS4EAmAoDOAlCZKwTGfpE1cJsHKFhrD5JNnJFaRCA00uaQBLJlO25dBahgwWtNLQK
2vQ/g7RYtugUJWayps26L51OEpui/OV6onkPjqTVI/XTQxeEllTo/xNKIYH+7qDXNBdrIlhA1LOt
GAxIJAt1yxoOWQa++3c/yUBZBpf4CQKJ9vYbeBvlPh4YV6SYK3wn4oPwp8K8TyXH1AcFRhP8A1Di
TfLSsdmhTrtDbNdWNmA0eW0casHSLSAY8Nwegsf5vtDc9OdORKIhr5hxsNAxEVIL32/rNaAlFZl6
zpf7IOKS2BHQiUWRgWEH/A9AlMiPIn4FsHtfSrY+/4JV0W+cK59rt6idCvc8HeweBe8dACAMZ3hz
lpCrm+goOZrZ9CXR+zgTQb8fOlmSPTY2+d9N4XDKcZj8PQ6FmyOaJrFPSlhSlIoQ2g7gdoWjG/wZ
7f7pEnvF781OD3Xy113Xj6TtRhnu6h9gGy10bxJ+7ghYXuEYwqNtlRtns9w3PZ4qcvvWZDXwDuSi
c7U2cz/J/7MG25I++rLvJbMjL1nVNfsxrhbukf4rYa9gZ/F5RuuNPQD1X/qdu1t08IJt6Ne7chQ9
/eKAnlDzvx7/zh2/Kj3kSESkG7AvepLruh7P2UyAooL+QxAr0Ajz4dVTnUnGKCIgpix9Nnz13Dme
yZ+1CzFFmAvoovQJIMB2QkpH6EZED7bPq2Bhf2az9GhlwIwcGOdGucBDmniQD1/WqHAmmR7eAHNb
7JQyoQPbAUvIx92aO8FnfKZUs5SF6HRv43HZvUXAPM1ZVukVMaAagE/jTYaUF0VVgYJchEY4g6z9
Ur2m9NY5JOMAhMxfAQsVU4kTSYQRlUrUIsdL+dnpPztYtOdwbNJPbStxPBikD9FMLPRd1tnkMDvn
jisuyXbUKRyLRoWxlkdM6RBU/VzgoBYiNvWo8d2e+OthmSPSqibtO3Fa/7RZ28KExDQsYFFJHLAJ
dMaj0SHunzzhFBQhubjj8SQOouqcZGJxXsRXnF3fWuqBSb3YgosHj3peGVvyNW6bgfIs6O37krv+
dE8vmsxNbLRixmBXqT82YInYPugpQjQf/vZCNCPeKYWiTmY6WNBHJeZTzUPxb4M/1YGzULf1hb50
oelKOErglzCOarLU5Hzo+fkibIvklvSBav1iiIEc4UP/okHmoUINIXCWayqUYKPdp0VOyWNT3Ei/
gE1PBoetcenSAcGsgF3qnIUejrsxPttK6vqDOlzArte610T1VMCvt6DDNQQAjkb1a8WGQzVKTk19
BMWXkOSQqyCpZXMo2VTT+I/KaiSPwnaYMB3AiRgpf4vC0cF9eWgGQHuFvDWCyXHIpqK1LsEQFb4T
FqR+5dY7kQQj/j9OT6pCJ2u0Kh5/1Y7pLF+nnSO0QT58P9cwuMq8pCfgmbCaO9HAcy6FLGbeVL+j
UZa60TCVr5ZYOznjpoKsBSQMd4dkwcyvWpLk/VGXIo69J9TPpG4zC7o43Zo3g7O4jNqKpaXj5FqM
QX0aTlZCeQT2addB3sJZ9KNDh+LOGm6hupl/ShvnGAdmnsKSLH/E3rwFWuNxLzV4nZ2zKuDseGP0
i0tBt77ck+MalfH1q2Om4ExGXrJGUdrleJrPTX1ImC8MCeDkFp8pFuKFoX64Kl4Ap6CBzrZjRK5z
wiR89M6T/cnb0zLhxb3rAz099eZh8UOOqc88/xUxGFzqyHtQKQvdnRaA7dq+GppHw9b9jeRD7+NW
0t8Rc8VrGH6ZzQWmta4JVbeJuYI0r87D3eyyNMuqVeIVS1VOQrcW4PYNPdQMVKj57MnMmNVEt9l1
Zhx2bcCHPx7AFZrt2WPUDkB6n/ZNyWiz3zUIYYfRtuI/jaFsdBO/iJ1E/fyGWWp1ZITNOGPiUh6+
tK5CETNgYwMtt4hp7NWEwvskl47qKgxSj07nGRG5w3yT68cW6x+6rL8TSnaf/Hi7aOtgNoxKhfgp
U2CH1It38pE7L7ikd0xL08AYzS5qlRdsU9D0Av7JAwzPr2uhW95BThiuHEfDXheVmN6SyFYVBktn
ZeUfBqK24F9JAhkTR3+7SEWTrQGZAyqvbojSCQS78z0pVHXEE+4ogHLZQM38Xb3x5qM0ntM42pRW
29Tfybs07ZHeB9cekFe7h3qrloycqS4K39NemuLG1YGQzJFxdJe8jaIhZLl13+L0AMBhjOP8RzYj
Xc+xhnq6St9UxqPcBpfh+UQ+pAgehCg+9jbgM3MhX99TIjl07qOwEvkR7f2CpMbh3HORLuLS/5ZY
C+LfTmwqWq00hqwhkhFrycdTjPwKmE9iOUaYbVO5l+PwE74TTVpHXlA4KHcRcydvgCBEYgnfby68
C1tk/GkE969zaRz0a0ztA1HO4CYFDKzZ1F4lQ0YsFVnjAts2NUT7SdI7ovUuEIto0ye4hxNyT532
n7MizOe5rWOStIuXCBpDEdgkZ7d6FKvTJRgoHYdQkZ3fvQszxEcqoN9WGJlMAqOtoogTxgT9Pn5v
JSSfSjK7trwe1+zHlP2U7xOOMQrnB4QFXKwAReEvHIYo9JXAt6ccXwXSGMLd8aNZ5Nvk/KfFgmV+
C5leK/yF1JARw+UHYqVuO57UrguJdNg829qyLZnMx++dp03/DIeMjwe+W+P9mYkX7jp4ovCd/glY
uAK1dicPj8dlYiy6bOBnnHWRI04NeNd1klw5iHc1upzfWDBbaV4WEQye2sWVUhx9M2qpnp1uwte6
iY5pqG689bf1tAysrrfi/fjtgq27eRYYiNc5M3IN2l9Jy1wfLyfDV5XwQpM6+6WYjOvtf3JK9Fwx
W7ZBvuuaZD/lRv2uf0kTy/t6gbQp8mhfMFZ1Lej2cFRqNQbR3+XwqgTHWt0xezFkpZscoT58J1JF
WA42ck2d/+6GNxOaR7FtggqMKrpSGYWgwNtK+iGfFBCjcXCJSiGRus10xCzdU3KDXJ6T7SOYr4we
cSI9Bd7iFbP3hyhwqWRrQrnWEZTdDOh8E0jdGEcAzz12tzosbkcgZyuMkErNYDxkXBhu6txN4zey
Opp5MeKDyhz1uKiFkjedCRf3pELDgQ8AOvPst+RSStWzwiB1eUYX3vX5chWlL0iNKnhJ/9JZB/AE
ZssOIN+NtDnMslKt8VFMDPJGb1P6FTqjQoHF1pe3k6Xe3zOgJBKfaJtNmtNWkaFSBS3ZORFBaaoz
NiXXUIunC0u7meTnFqN9uXRCT7bVoxSaZk4P5oHanUs2t4YXMFFDyLQWM149lEr5U7loXPCuQRv3
nGMm3SE6ezNtAcec/qeD3ae8FeqzmNGI+k4Ib4lkNBHVs7+L6MMLLYoOiThlKJqJosKRi0KEBwHf
WAl51tnlh69Hk0anQhKJ5dRCt1nRJJdQNkdJ2/JraK68fIetyhtl5QvP1wUDngLti+H4pkxeHBZA
kYqnLHGMPgZv7OBQ3KCoZrSV7TLaAlMGN0Zy3f/WTUnQyny6a9XgERuQbyXniq221oqAI8lkUR/6
NCdgzx87C+dUAL5IIboqoVVWAKKyv0pggPkRlPomdQsPTg618I4pb0ZSS/G/1h1sYATb7qmnYyfR
st+0GN1PIwYvROw59H2v+uRI1iR165RJNPxNOWvte95v3/xBgmyOKPna+80RFhFGYIeVCcbd5hyk
6moFfg6HKsQRP+oERW+dOTzUNXjlQ3JGq1iD8S3LqLjmT2w/PnM+ObeYXlMDh7VSIZPMsKVPBUiy
Ry+zlM+R7CJP7aV2ShC8YmqVSBEbLbWWufKXX3KvUAoWSuRXI4qGFueVCSjjs6KnwXBz7WvAHhQG
v4XvzOfp8oiwC9yc3WUs3f+M61JOh+jNQkJZv9MO2QgSsNxrkwofmIs4GSi4BjeCurXn1z9DyYu1
LWPsXWRXvDiNawigt85JkqZBtixDj/b3tAuf3+C3Tbafca+eMS2hDBHZ9Q9WZZNsM9a/QJQQuQaS
8RNn5PhfXbPMd9iwKyyrGL0fj2OQVEqOKmK4ENyWVuYwv3JlRYr39WKqEhgTQa7DZTfQCX7JW/Wi
kIBao3AoqLBZBiAZfFKaZmKVU/cjBAuaOm0yL3fQ97zYnSL54Djuu74PiQf/iDR4/Aywkots7y60
lRiA3hfyF2OCA1Mi0B7sEJjm/wZJNC98Ejixss/vj0TxKvhR2Y2FEZFOWtOH9cv9pd7t7x9ctwqg
CapTEpWYRop8RytVNXrZGM6hvcFIE6uKqrUxvQDv/FgE/2kdMhZFD7LowOAAOxT52piPhV7jE1ba
5kAXsuOn+zMeMXdwFv5TwU4jMGkpxO2WSd0JPinpYweQp8YJHiG1uj9RCl3hcV8ArAxlRMpDNcxg
GddyqOf6fcXVVsx+ME8RXj5o50IMLjVfb/nX2dzZ9W7uNEWlsHEGHktacqyvTg8BTZdkfZpjm9kg
Dj0DW1/N0ubMA8SqrdOUTyh8k5natx4jdEZ8U23Hw655ajTnZtkifD1JgcVeRvJ5pFHVVK+qd0MU
DT4slh/Zz5VVpA0RQ+qvW1zeDugWxLPfnL9MtTDl6sDp4LSXl+mAKwmcXPQ/vqSDthOut/+g273S
KfYI1Xbibiv3g2nR1+6YOd+8R2+01+OwfboqR9XO2VrpOL74bdpGx/rKiKSrePedCElT5Ji8R0nW
+tDANEmlQek3l6dH+On+exPHvr8ILg4YufPGRLJK1Ie2QwOMufbw0mDD29wNfdctPGT+3qipF+5o
vWnWKL5YhcS/4F0FIdci9nEpTO3nz/LawHoevK6kR9nIjsBTB0Y3JJe8p5zgcVdboock3CEAltIu
C7SrMS4skzflqCYyoCadrzDbeFq50proCzdxMaFSzPIkipPIS1CyJ9JNhSGKT0J/4njGRwrr0rlZ
fzXe9pS7zLBQU87v6ks9lDA+A/RUHWXYvzZKFRAqW9bUKbhPpaHC2qbK3hZT3aTu6r3c/ljaGOzV
TqklQzRMV7Jizg50xPZRiciwN42SVKo1NPxy1nScEXH/en11yV9xz2o8yx0qVXEetmHa+2rzp5J2
MdsBP/bZOTyB0tdhKyU1/8bR0tbEyFJil6uuSX9xgfP7EYhBu24OG9YBvJ7YS0iU++eK76bbMTdP
zH8UhLG+XBsyBZSFsiqzAeG52UIiRThSGYBioDRt25VwuTi87BETzgs4iL7XvwUMj+OJ9H8+SilU
sW4u/vkenVm3+zzhOlZXyry/OK7+ojOWDoqW7N+Y3m2ba42MEiWL92CYM0u+TaTnP4vMw6U7YHRz
S4i+YdogYe89510bakpJlQukhQ9BxRAYw+mqld1I3pYEfmIIlzpWTrAnUD7ZJC1otsglY5b3e8cF
XsGNypNIIa1z/cc/goYO8pJCCqdG+WKDiOM9Him3De92poVqTH/Y6vXDdytGQnwTziQbrG+U5D4R
yMMlQ2SEyex0Sdo4FcQ4jpOGG1eCyNe5vOeNOh5eDKeqc42p3lw1egH+BvIcgSR2+g/c6656a2hC
YBi/2mC4cM9VhfLvGpkU0cp5cb8DEKv2WJHYojS+31/DGQL2qehSJH6zmO9qehfkMxCOZhO80EVQ
EaChH3d+4zV1jhieoxpdsptf3J8vdcRFtp9H2J+TsScMEQlOhhjjgV2mNZI/xSb35Cro0UPIumZS
XRzUHU29Sxgi4lOB+IJbH5rHieKDU8erSppgPdAD1ZUtEHIZvvWYpLZnhezogakPxzg/A/09MtUf
Dkc3gn08dn7vby1U4LCXI4BVbybWvArPinFx9OYa9Q7QvgN04Ws0lbEn7kIXv2re+bSoTFSJp36e
kZ5pVmonllUa+O9yWS8LSNS/v6d9WmxRypWL/RvOC5A6pxOZO/QU05PQkOpC+uTzEvi+eN3vK8MN
6R+W/TdtUW5OG9zfF5c4w5pZUxBdwZBYkCV2yBgx/YDbQT6rl0d35oac34YXwhNAbrv1mDk/zm6j
oWYJrU6PSDNPzlLROBhJxqb2j4Rqp8EIoNCqeTU8cw+qtk2/sSowWw+U995+Iq/IdfPzPY8Ecf+z
1wKTSMsEM3ozqZW3pZ9kunuM6BhvGBpJISJ/lcJZDy/TbQOlkmJANEp9cdyJAnbQ2FfNXkDZPQev
U7JewgMhz5DmmGYrabdNBIfETKary5XZvWL3W7Z99+T7+t+DMriWVuVHWNMCtMBzoSxxZ/bQVglF
cq6HfKYJEOCV8WOjB1jyxPgg8N2beScGfSzyMm365hwcpZozk0ORIqhIrwH9iOwx2QiwWh2/zvPS
KlAKv4E9eI47DIB63sgnWVTc3D1XnIT5Xxoiouzc8jry+f1vxOlmNuc2TVCWo14uLqdmWOSauoLd
S6XLT3LamDRtEQhPBuw94y/JShCbk2tmPVC8WTRd0LiWJtpTMDvtyeWrO3TM1WiAZvKQ2KhHwCpi
oonTDqwYHA+dnvCC0cAQpc/XDlQUk7BUD6H9OYFNNzcpwzj/5DHKgQnR7iepY3ixv1vgXSRORGvQ
hjBR2pJLznuk2Wi3hVmBXrpRj2HBWV96hm3Wn/25Roqp9WrCPD9dt7POvs6WRBy/zBO/GGX9cLWc
Or9tJNYfMBBNLUo3EVDu/sC3T+qylsILjH4/qwv+zZyyKbQMzyC9JbtfLOAarGjgtOa6K00bFrwC
BnX60OBKrXsujFDGP8lMEv84wPlKUOaBLGldpYDBEvigNt33IzNlnmks1jjKMhtgJV4Gyv0fiDio
iC1QarAK9g9emrRkvH2Q9DrTbDuAZ3i/NHAsLQfsdfXf+YzlQ4T2fL9mJLEKL0maly/nkTTrCY/u
XOMtZuRPjMpVTa32ZmMMMgsnrQqr9fPGd2TkVvgwBe8Au5E7t5azNgKgE5ZWbMZ5zHELJ39b+0+Q
BMSw8roc2M2guhE2/xJonr7cUaiU/hCgPTl4GPPYqGNtlVTsvQKKkT2zmxscXK21DH9v8Q6u9TcB
WYW9+Qo5nHGeK5djRN/49HO2a81HHhLdezPdHe022y22Xapate24YybjVnGdXEIAH/Hi/BjhPDXc
nC0828RMlb3fpgXojm2h1lhSKcIcIcegPN9XD4SkDj8lmSDVhXg+/aaklqWSmI2NADovHLSm+c/P
JGMjVG/s1xcysc2Kxor7hcSySV+ZbpoaUHYbFxBZ+VehmNSE4Br3McYzcOZXdol9pKSsLVyIg3+h
Yoe9jw2oqPegAiiuU+uggIpiHgmPQzR0RMO17v5bIzD5E5pDAOhAwTOyWMe4RWfwMi/zheTdd05H
HgC4SNs/EMRZojKOtz5KrJ/mpq56FKV0Sh0+Hao5z//5YS7MWS4GSXtSzEUs2ZHAneDsosvZUoYF
2KM3tsQC5yzmQCF0vnRCh9e0QnTJM56Z6KhPsNmb5hs81A4j18o11V11n0KmEFo+G7Qh2XnGPcxQ
4Mbne4nga+jmNyDKuvojtDJmT8aaCCwwbCCzNR7hSbm1hXjBuAuENZI/W8tkhN/tlSKjAaB2EYNN
AVBwlCNWRskQIbVLZP6jBPjvNwIUMoxBD4hh1R2rDuk5V1MDQzs+PSDXkV883Ah+HtYDf/tvdjnB
E+52e22GFkBzGyyRsKBVyGd4Ljksn2kpPOC3Al5C+5nV2ApVu2bP70LwZ7y5ShFUBoFlTBMEdvL7
X55LMdZtNAA5NAnMzaDkP1Qpwt5B1F6OdiGCqGu/RIdDGYP5k3V0fsVrkdItWYfO2xvU9y1KeTKi
p3chTy6FfDREYl4+4xpGCzeemxUb6wkGjYjg/UdoTm0NtoAOTJao8J0SaNyReZHRL/yfdQGitBq4
oaGacpO9cS6vhQYGI8HXccOdbPz6Hf2q1bb9Cux0PoYpFqngUUiDDKrN3IFIRZlgGLozpeTr1k3q
n1BrQJnYsi1S+P8HHTzf4GducjkaVR0Lb/zM9EbfFvy11KbLCCeaDXkVLF2hYtAsw8zHbtbGinVa
UpmGyAVmAc+NQRfNksep459gypezPGjxBQAHw7HTxaELIpoMoBAXvbYLZCniGzSfUWMV15mZkFVw
xirD7RdQv2XXz19kE09TtriN5R+nQ02NJouyLpVlGpkaWK1LPBgvX9h36EkGADuSo3WhP1gInZPC
Iddu0qpdfhUvE/2VxdXPmkVazHUcFd8m92h8rQZibmhnqOty8JftvpNlzrdt6aePfG+4O1RbJji6
iYoQcdfzMHnFlN0QjdldtJ3P/OUhMgPsgDfmRKqKfGw232+rfz6OChuQD+IPqJenD/HiHm0IAmzi
5x0G+ZACZjO3q1zLIqONEgciy8CCCf8CgCiu536ho9XCqUUhFQ0cnjudA3ngt1k7WgXPJ1v1RtSj
+/cDhWs/GE22p1E7YDH2g8YnOoz2YcB1l5Szr9z9NeJAxaUForcVN03PK7ONVMzSIyKUbVd/SGbh
0FGJ56w4ZC/Kk3S+bXyY7Vnz8syjyRR+jkhfAUOz7nMfwf8hgKLXeVBIblmLowpjKuaHbanOw3hh
Uy/NnJfn3e4QRKGuev4QKKUfncsJTq4AlqjZySLvUiiJ4bxQZhKadwRGLM2m2nUGtgxXjEPa1wSq
ph37KpiQj6x2fiqH1oChXvvwc4QNhyCeXiYm3gICfkWd9cPHopqZfgOxTiOKvWLc7llskAK+TwtX
7jUIAMNAjDo0MnFwSeRuMSpsPoUPUW4p5pcy+9IEad8BzDcARsNXmVfdOy6tkcOpFyE9RPWtxElW
LWw3r+pi5au85w5cYXvBCU/pGKAhfgpw66oa6WtBVJrwGDioGOntr+Ut5HW3tjD6sDWDDD9V/Vym
S3qgzuP1F4cjppeA5+tpg1B6vEumiYLfnnjl6swqthFiTI9DFsvYE7oSIuMdmfOwnzDdABIRwhIm
7KT3yfBsIJDqT911d0RoXCWnQEJD1KpDG0R5BG6hikutWrHudw5Z+bA+9CW8oeEOC02hd+ZimPpO
Dmt5Nqo3Km+BjSJ5eJ5mS5Prxd6eh4yM7+5hIPz6yDTqxSZuzlzIlfsn+ssgdTCNWdT1GNYJunWF
KrdFmW+npELFGb30n6XdhIcXiqyYfZ0Fqqsk//OS+f2qc6EKnszA62ii3EVVPOoers99CF2/wEvQ
go9iktMMk7srhR+sWtul8YZ7jXDBzPiimSUl8YD1dYEcRFZkZ5AyKYueq8HHrRN2ZagZn3+rscDZ
Q1mJ9vEnSWSNdFRla5U6TbnodomMKv45MRQMPWiOWJ5+f7t77ASXW2D+59dhIxWjClAYVg3xloG5
9ZvbLesF9NYp2XwD6LiipK6Ro0w5qd+kTkEgXp+dQ5bJi+n25wTZGoOGo5GhmXzlOAUv6JT1Z6tx
99NZEzRLvZV3WB59e3koCimi5iftD82q3B0uDLgZNY9LI0KTpFKvd2r4vh89LDKq4kncKUeObiyL
Tx/nLWo1UJwq/5Ir2zDnmIcVhGJPtzn3FJSO3Fj0WQMinNooMLDTBNTFKHmGGf/9+fsayN+SNh1q
URSiFrcDq/df9PnyEofS0wZ0zgJSilGHfGdLquhYcxja+fgYYTn8EOTbyF7DWr/gyqHHmENcHKr+
unSL4jymViaALrk7Fsq7fHNjvjtLF4OiQxKjD3d6uE0kAvf7SqAqIaey0AGsmP5IpcvXe2xii3FR
/JkJ4QI5pz8owCQ5jLgedDRLQiJUnYUDczOLljhSJzWObbA/oUvZN5Mf8ScNMmrgivWlgTCtuQ7f
iToJKvFGTrgZkLg6/T8NeKFGBfjTLpqN6oVouf5mtq+0At+t8l1/ejCzjBJ+elz9wyQAe/2Uicfr
S82kBOEkdHS76jFfA878wi+FOalJo10PJH/e8gJrGNfloehWgyJQdGroB+jyX4+2hSuPel0xWzB0
o/FSD1/IIT/8Q+AVvTb9Q+bkKjEFpAGC3/J942uYjTABIlAUysxKn5JXPPFbbIY0ji++GwjEHMAU
HJnr1SrkdGrEFiyVkv/f++laH+hWWfhYUFLIdeBp9WykBP0ngXNjTIG11Fzgw1rEH5/N9rjlPHlh
0YqVQlThd0iUq8fgx2QhwZyawnnb2VVZb+cIwO92DHxou1oq116tQcUjmLJOg1assDwKR5afYx/N
B08DfJ92x6Gwxa7vYy3LhRkJs18masVY+cM5cCzU82WYa8Ruv9qdiVdoZs65MP4F+RhZmEYi9atK
UkohHDat6EJ4Ikqy51tbglGt6wISddpsAQepH8Nxnab54sYDF8pdHroJL3rwqsyVxHc/iSgu7OJ1
8ixvYcx//THeNXjO3T5osqTf0KXLsf9oviBSnFdViOmcxsZhauvMcgvNqtKEy3xeWDSnH3ajkm+d
CLD2SQQ1B+NtRkqf2wJNxAQAe2B5LXASfdhYx70qlZlbkBQFZ+4Kp1w/LoXLXYX44K3RMixj6ncf
heIKIx8CgmgWGNP4demuaz1rC1OQ5IxPjqU4VQjmxDzAeebDLQRvQR+1T/KX1huw6S4Mys1H8VuR
LVllMjwMFsk8eoEICHcKrmsh6lp8JY7Leeb9kdqakLatAP8cqgI5fO3PNcOT1h+IDVjr77h6kKdM
NqucoHn/lNwa3Ghxe/3WssKNnS6Pawm2L4qsu/Pw3QnHaHnrdt1aQYxcY1gZMUg0Im0Pyqy96Zto
6Wg+V9xgyhnJo+GRK3wneeEekvasJgLb9zXBxGVWFA55LqLTX0nX/jUfVKNGnBrwOR2TiNqCBFbG
d/Pa40Sx7SxFiIiISSRcK5+Kzn+ZVE1i/5gcZcDiiYTSJyyrDxe9MPIO759+FJteZy6m5KxsFKp9
LWoOPimFguEE6d0mCzFdPvL+9/YaeNYwKAvgGQAr0Me9yZhgyPw8rrT8rFwDtFJtqefRfdJMt+x2
grAoByJoTJIDz1M3gGPxpa0zH24aos8iqW6U2zVlSgKQQwqHHG10WoOBMxG3rteFboOCLz2Q8Jv7
3TSpNU86i8GsES+ylP7KXsa5dPRZO8WRjjh8eTnAOOUg7YbmWEp2dhLIIrirebKak782Q+kmZdr6
OoE6nLKmOxC4e4NUy/BZ3KOAlFVSZUl7HJXgUo9qGfHpHSn+lODp3Xrou2F1IqZgAgWvlMR3MJf5
zqjQCeQEJfeCmLCY/Bb8hhMiQCP/MbHOwdH9Q/7HgiZjHbnO6PHKuLkbjoGetrsszyCvN9Hvlwrf
B2HohJEdFMKI4bCpNlQFYI5cbwNkEbc8gKbifAfBES0hfotdrzQc1MqM2qBF5L4MEwJrJvAaSEYx
UBz7igv3ZsKmowdGzlHjz6mU8bOxLu8DjyqZYabGJrORDeer1d4EQMhr80A2Gz3Wn5CHNu/6sJm3
dKXbcwKKqirB0jMBxBANsJVvvOSny8Oo1lguZq55s9caCZv8t720M3sknuBmcYz0rezsG5aJ13ht
IG2cQeO6vUOZRtY6ikNC8Ngzw6tX+T20IVGWX7JPHh6ZKS+Sd2xYDQa77QhweWLp6nNeb+coNPjg
FXQB9p4DSGnBYFV7la6yXcPvM1nVcLA0Fn8aNy3fRQpDpWPYCr2CgzH1vDSEBqh9fQKFPRER63Fj
s+SdmSNt0VUr+3FGRuTkz9JQAcf/FxFHRmX15Bdhmgmhkh49u7/7STkBaMEhPQoOIK8jjSDcvuSh
nf5pUmXSbLy6fawJ10UVyi9jZ+Gbf78pNV6jda25ZmOewut+11fME+7muJhg7rSN6Lk7c6MAU8ir
PxGbnfh5nUGOflZK1r9BRgnpado77Q7cGmtdnfIkNabOrispi7KfwJKCuyfv6dyxGDvfexgarzNr
Ijhe4W/XL2Avc2r7BNTO2ttKXEPsr2dSexnETVXaEpHkTTJa71GaDQH8tZaOUxLTDRffHjZVnO7/
k9kLswvKQj/CayXSh3pxvboxYoWSH5tG/ocijbpMAKPQTpCCD0jL6Z1pKTj+10PHuFnb+Bgq1Vsw
L1vGVLWq28i2SUyNwdasV+YTG2ke+M9zWfVFT0vYbLNH5O5GZq8en9TI9qMAuazjJyfReMuJ3IXw
VYDjw9xTPTCEkefkyvKZVuMXnIfAqdfCb7tJJ/YzpSaNmDVhzYH7a7hPel+nTANDPCvnhL7XJ6c5
SPIrh52c9nTVq/k7ynv/4HlsRgDgLKFPMKhNLTGCAFeJjcZhGfAmpNtY+VOvp9+2g/Mimw01UuHY
jPgxlEZX0ZBo23RXgdmn46gtKdWPFVQnj/kCXdkTbhUsSsyXBuhwHjyy1vwtbeduf6BnLcpuP1Tv
d4WU5RcfnANwNGtqC6m5QFRuCGhW6seM5S7T5xNqGMkV2mNTLRejXexFqdrKkbbda9ou+78GkPMX
KZSNrE+P1KNqOkDbEvD5dYc2tjW6baYYzlbS+eAesfxqeL5/lw3ebnd4ulD0435tz3Pd1PXvezCh
+AHyqO85Eu/dnjFPNEg4dO3AmLqtVZPf0JKCjCEUbCHPzc7P62JPtbaTelyTM73Q4Wqe+Zf6loyQ
sjhGW+FLG0skn8CAsGo2C9iEpeVWoG/40yMvKG8j9CSo5NEunm/XVDdAX1LlXW0WP9ntreiOCnxA
BhAD/wtgECUfNI33raaxA+dIL2Ri2U22O+sfZUR4xElKwWAIvHUNoIIw5WlSxX5Vwc3wvuqNZjYq
HkkI5yMeGtdnEwdjLfpCEIgJa7S13ccuT+5dXfXFC6Yyks9C4KMD1sJI+CgTxCJlNPjZmNHWbFbU
IJ783v+rtBySTwdYwWQL8Bre8lqdzVNucMJI7EOcvwXd+uSFiwwyVs38dNzXWAPykcjqSQb10Lg+
JFQqzGr5g0cgg9yFPrOJvR/jiQPl8STNI3DmCzvEv4jR9bQPV5ozL6Q3OzIACqxglaO3rVlIUoVA
Sdr2xsJRr/3JEUY9pecRBgFRJfy+V3aYouyCbEo7nrX0S8TvVYKF8WHz/QnUGK3//tgiggDiY9s1
9YU0vbU8R8SMe4jSZ3P3kAc8mi7DTUtWPpQH6XLS0W+fqpcPIc85pxeIwb8wsBetuoVReRa1SUDZ
TNuZarpkvZy84dTLiPyUV3G2ujablxoakSNUuEBRu3nAhy5aSQK5oarslJwCifmQJyVpO6/jayIb
SCFvnlz27bab65Y4ycC+JBH/BjWcxHBW5fuEaYTob6D87V7aF5ftCVObaf/zjG+MJp87Qpa/YXpC
AuglqUWEz9hl4ZGoiBA4x3q4Ni7XSPqR3DdTWa152znPzGQkYlIhagnXpM/ljKi/ExmPrkZPlY6t
bbTlL7A/Rtyxn9TivW0sejomF6dTOz8CH3sYsQogJhr62RozMvq68VMMxUw0qvGq5Cec91QBcL3r
6+5SEsSy36PD1QOXOVRR/EZZX112fmLn+8BG7PfMlwTMrFfmefmqqXPBQ9hxv8wmpdqbZVMq1Dsd
w2n6ygnEjFiQn6StVhFIGUyvZapQ8/hkgaeJ1nbKFl6dyFEc4Wt8RJTOpyLYz3c+2Ce7YHQyFOKO
4JW/QGWX202AVK8NpizJ/B+cNbQb6ge2JicYC+IY6LrlkhS6O1jz+edrBoh8xmypnPZucVygKiZ/
Nnjbo/xB1GX4vqmjJ/LuI7dwWSZP3gz3S85IcAjkI4zxiszkffq/icv4qENDaWZ1E3lebLism+Fk
K5N2iqHw3Nk8cFa8hLh80hoZI5LOeb3eRBaSMGokDL0ueXebyIg1D8YTAWfPjR/83u2ZAnpcxeud
+9dnuv6CoL1UZm8NqOL4uco6l1d6it8LhQR0xOnYuwSKTi/kcKQkhdncxuvEnXJMC/kI5VzPBTDD
ugnWz/uYGlvgbkrcFkwA9XGplREuOABTOnRuHsu7bMDxbxOhG9pEUElyk6BE5Qn7CiGdht8VGdAk
mRkzZShhEHHcKjoSug/71gpJ81tlshwqs+4V3j+vYInxBkCj+C8bTbZZg5W3h/AwKTRfskjd3xs5
gRoGBRZqSsSXzQcej7DrzaY9N5RIh9W9CLJEnqPlaLQ79XYa/fL4Ewzt5tgwBaMe/JLjIHl79pn5
EHHqP4s3pT4UsBtIIYO7On2TEc1r+QvwDEo8x9Jz6LG8OBA2kohH0CCcoKR8ygrnDXk6Myw13Vfa
85cI6SEmOSaExifuSPxEtdTa0ro3EEx+wUiReVFlEQSE6BLb8zJE23Gsx2N9b4J4RorwGR77Tf70
XVHDy9BNPlhRBAgYeJaz1vZnfG1EnoNo3aG/gpIW1K+OQidy8cAjr0qQZLzrbmbMEs/atZQRjtUV
Em3cPWZ54zdJJZgcBYxfEdznxwu+NmN4LWWtXOuciI3m8fDmCcXoAvS6KPHIvSo1LjWLS8pwX0nV
yTpVmzB/wPWCeIW6Hq1SpFmw26xvFh8DcA8gehSzeB7R0WTGEXfzYN4OUJKdZ8j18AGxcVHHFC1U
hJFhHswJAHvGOaBNAK+efjEF5KdYCr2EnJRsTqyuXvxHBzCF6WJ9SIQ42EYFbYRmG+iLNjifKqNI
+X+Z6iQZna4hyTId7Zp8OyjtlKfIZWg8Bc/K6jk9fed9z0R6cSgQP+FLNTgp4Nin3GJwSUhu+vrA
2HMlBUZykcL0o0Nuw/XSK4agrfxL+pM8LGJoQnqaxVgeAzppM2fCFX/u7qBxA/DztNFId2OqjA/o
06iKgEKhA68wzFUYa56Qs7G/2nrjl3HQJ0XQ4yFP3LY7bXEHIERUC4LIH4bzgH89l99MdvXEYQa0
NEvXm7zDCqaFFiOJiCyuUiHGhBVaXEKyt7vaIcEZbVnrHclAUh3I8nNmXSjDUu8pHrgR6+iSIvIB
p6T9ARWZngqksHX29sNM3lR6Xgrjvi2OtZUyKgrsTAgM4LcYFBPCZYhRtxE6HD171X7LSUetXEB9
QvtYwiCk6rXdpPotG0PV3dpBioVZoLudG7YMX2PdUnQE8Zh84NiD2t6AUP9QdnncYG/b4guWAvT4
LtkuaVlyvuvbb1tt+DAjL7trUBAA4UsWfm/qp4xJnnyGwsBySxw0OZ6n5/qS+seNB4GWinNO0UEP
/43sMWTJZd4zmOPgH8PuO76bNfJeYiVSsQy5By6lUdRmlgS3UIKov8kPuGkUhq+6ETfBMG+Lr82r
abO7kcT7d9/NhizpzgfqeNMlCNzSunNLvqsFXcYuRaXyzaQ/H+alZ21wEJsdBp+Uqb0oC1upBcb+
mela2gWsP5jv7W/IUoPKOjQv8nsBhk9a9ykQs8m8PIYMdWU6OFfbTJwqd5xmGfvp4eGG4Dzy7YHj
KrXrFFSa9KP3Fj5Cnvsv/RukhdWM2ITs5GJ7YiSlqDJklZHI51pNzNuPZCBkxFe4Is92DhI8zGj9
gBaFxI8XKZDrKMve2vxDXuPs8TjJlu6/7aaub8k62Sf0tar4oEQrquLlwTGmDpoptJ15zDwqYEDE
RFZk5mVlf9wROAA/to2DeICdf9BbRsrz9vRJ+o2ctoUJRaEx4oAmjQjwRkxqIZ8o1+5GZ7zE8eVO
04DOv2d0Oktl2duzy5NwXviNX2XnlQBY283FlTcfnR1V7EvOSdeQzoP3lYb565tdIrztjpktx/ui
bwBdtSDpzrD3Nb/WCYuIc/xLnC4jAT4yKiltXk5G8DUpuUqxPKm0BL32iHXo8AHgWDxeChiMu80f
0lmyhKm5wWqg797w6Ktk60F2oG3eWk/Kf2gZtu7rTETJ4qaIzv1zVZASUZTajbnR6mkgpcT0NMbU
z8njQ4lK+7Ha6PW9ZomMMYddzZ8uzdXIqqu1nk9Xu8sc2+TRh9/w440spxocb5GdClUzHKVDPbb9
DVhmy/QfSI4U0wxrfY05a6Dh4Gh1i+349GnNICN+ASsAhoNWjBJFLv3q9Bdd29n5G1XLDBMee3cu
FL4NTjqqM3FZXJDZqmH7JPEO8ws9WPQvi86xgCYOs05/GGWUTj91OJrgvfQpXw94x083lJOvEd+G
wmTrrJ3WK5bXTI/X3/o5oMuDFqGpjkXy9i+itJYsKWE0qjNsDW+Ms4GAKB8K3UCOd99y35LWBZt8
+6L4jcrPWYW5Y24yepwitbGydzGufbSDLCu1CtmvUCpFzOFO9TfoFvW+Z0Gk0aCotBGzfOQ4t4h4
3LMZ2gxOlpOI1YF7HrYGxk3fhafElCR3dJAa0p5fZlynHQ2H1KTvSINMO8mNsQ+N/qkPIe2ki/6s
ynqGKdopUWseUANzHr3sCMbUNT0lf47JlP+cXhK2SzzSRuTz0F0U4RZ0aqDRNO9k6Clckg07slav
zZDqYyCIaXCTLvp4bip2+PUhBA/Ln7yzgOySM5lr8nJkCIjkusrmUcFRGkh5TibK7nUZ6c+7p5+D
tZwnME6K2nfs2Tv3uIds9w7zWLe1bubx0p7QfN4dXkdDNEl6ft/O+M/vnVIx5mn7k8wsBOK8RDtF
eoExhvwJ17RG30t8vWhEz8qBsYoiJWwPAw3+pkFl5eDw9E3i6a0COJTQEBpvhDRmKn0ArRdU1taV
B2Um9vihTSGxpjuRDzHyVMr/sFuMxWBHn2GWLwwUZX7zMaYebcZIb9CE/Rq7jYAB/wq2uujtqLV1
c90uZ/Cqae620Pwdwr6e5rlnHaPzvdSR/FfHNtUKhxuo9ppP/g01lbWcz2q9GVN+ShEXt/fZs29W
7f88ruZNWb57hJlNUcLuRPGaTFZhs+JQQH0vx6v6juGN1BnWsfPisYeWhHt9oxRZNHwiI4jvE3g9
MpECh0fVLgxXof/w0gN5Vvz9DGlt1gSjqmUOIRBfhhuGZ02sxCKYHWP8HzgpUflQMvLQj0XzQCcA
RX+UqDDUGCQpfCQyFlZrKm10H9gZIfa2D0tYNfOv1Mla8S2WWIkyEjOYRcBQ12w0U9UAb/jyjQUo
+7W8WnBQ0POU+f7OAIztLc7nnU5mJQTKJoqQ2v+nOBhvYKFEM5NnC/fEMlGYFsnGR4kqjmfJ+3J8
BeoxOcz7uedSeg15er/Q9sqzZCnrqcs90C/8UakRi5Ryxj/Wts89ahor2etaPBtMx/rEf904auLt
LnIceYnF2h3TfWhZGDhrZImQCRXG1BwFbmpqQa8dqX48lVyajkwMdt9twnf1bkDWZpqPcE+L4NNl
XN7jjRbLlHA8wRgsd9LRJHFHkgsznxkwWGzVj+xX2mnz6bs5MgbtgCDMJAOtHxzft/lOyfHgloPg
PkH8GDU4rFCs+ICD4ML1+M8rt4XZMcLVjNyrzL5kHatidJNWObnF4YzwmwkF0nzj+Cgg7m4kqIyJ
Qr3ZLIzh/KEvOdHg0Pg+BIuCgwitW/YwZzaVy8mAEeE4ULpDoXgEZ/67jYGEZuWKfVPkqNtHCg/5
8+vslepg+o2juY7KroMJdbk40Vf22Q9Cz/0/B1sV+bMDjipqiEUCzgPOHLcJ1fSPzbruKVYjJh1w
X3Li72OQIx3kSKFsptcSt+z4Grl5l3y/iOYa4xerpfP5olla8NvwCVhWUTiZUf/Lq9A2yZEcYvPh
9Zcgi9MitR9lacjcWxSxnmsjV6UvRk6KDPUkK2puDuvpOqKRAPApIdiHWwyd2WdpFAlt29MmpdHW
oEFhxSEX4jIGnmI2SomvImExhqZeoG4HheS1V5iFDx7W7g50msuMU6tpkxSc0gTQZPITdgwg0/Dy
EmeizMX8PV+o5+lTvpv9/9RAM7DOY8jufZVNzJfZ5BptE8OQXe9hcwQaeTiZmo38n+CsSt7ZpQxy
XSz7681tnH2Qqi26iEmxW75/Cb6xe+rf56MIMfmPE7+sek6fcd3jhIYnasRd+jrerjiuZDgwnJiU
jL+OVDtwzIVb7c/qHvSjt+/JNwlpFJBBqipDLX+aWR/tzQYJ9naeeTF26HPpeUKpKktfRiHT4ZOR
c63tYSp9m2CQpqnlflL7Oy4RDTGuSX4mXkvqxxL7UOHywmWC2InV6jCZ37TuWXfiGFWgOPsjWRf9
y8XM36616JsJA3dWrNx1ME8GXdWLV0Xt7utUsMjcQEEAVxuiZa754XhZRm5VV9rz9zBb9HGT0pdF
i03RdMFctX/j3t4cpQppqVit4u4pLSd/KgrfDa5te+n8mRfP9vOuXw8N8A1L8AkSHC52W2yEBCyR
1Al7gpJ10xSFXBLtyTeasPJOTpuTqfBM+HFnuJAUbuKaJWaR3VYEwinrs8zGx0JKBVd8T4rs8gtH
uvmnZoy7MauzxwkXv39jee4kiLCL6MJ65OVYInLvycLKFjMt5N9HcCf7G/AhFnuFzakhg1viC9W4
tMiaxtuRZnRuQmPvc7ghUXipzr5eQNrppgL85xdZUXg5H7ENORE4fADUGEzvy8LsMbEs0ql8KAhU
WmEeMaMnNQAc7AZ/cCkSSAdJePgjAaDXoY00IH2bVtlaAgLUEufkhIRPL1oK3Wdv/huB07bb1MFz
VIC+sYbEMj1caJhy15XrjHAUKvgWojqbHkJJSawR7+1DS4v7bxexbP+FEgjv5FI5xmd7VQtHlU0M
a0yZ+2BDaEZKDXLTeW0HKGYUJ++LdOrHcjuQL191b9rhTGVaiioE7U6nlYSz9d6q0E3luPpLmyi/
cn7Geo6/QnIN+qszWzpnS14C6T0iH3Xi0ya8J22/01EmH+6OuNwgtBDcMM0q/NzzzVtd003tx5pf
ebaShvXubE+UVfThPclYKvSNmNTJp4V4FI1HZudln4LRL+R1k/Xox2zKeMf0nfsanQcuAHvAL9Yn
h5b/Ve8YNbD0HAVjGu3fPeEoN7xCYlFbAmX0RdVVI/zH7d5eWolkaLfRbUQGdjYWlbZUXtUTjRCU
SY0SdhKbdgRuSNthvZjfQ1pXebf5NvH1aK3dkU1QlrpvQ/5kJbAmZxvJaaGy4v/ZR/y5y+vA/uLR
EMSr/rdCzxjuz3gB3D9L3s553+dZes/O7VeeZvsMxHjPe5pOXs83UQ/mUHX4mKlMD4g4LhqTX7Aj
UAmXdP3GMd0uffbbEa7SHE5YNzu663QW0NTXHDRtmJxPRbTcBCTysLPr6L1Vkp9VRi0zY1MZzUKt
u/w1Oox7h+lp9RObfCsFhwvn6MnQTYLCRGbbR5rRuj9woNDhnnLEV7pU6PoMT4fWVOwKhxhBi6Yp
OG2z3W1khw86wt6O+FYi2EwDAFxzD6JlZ5NjR4z730jseHpCuXebh/+eYBW7xWmvlp0yPsoQPNHJ
2mKKHBpOlyM1Hf7kqwBM3eXg7FkswUd0I0yg8FLB/wUWD4XeiqJq8GdTZNIwTq2oRZSwM3WiXDYc
73Ix7jpxKGtHUSf6FYRU3rBtn1/NnQKI/MQiGTbRvptTpg6TSwXMIP4+KHqJ4Y6hHLtvRyTVLVd4
kbN9FFPu9T9ThQ6snjx8VJWV253CUDyhVHfi7EpSc+mgn4MuTlee61TkLqA+lT5N2fx6S+1NWmcV
5UAeUrmZ+q1w0/gh31OFl7qY6/qN3AcZYRb1ZhpNuYPDA73KafVx2nKB9jOD8ET6CmGYQ6kCCU5k
cDrW9QeWPSLxphC5RJCGgMpBizlHq3G2W3n/B1rDL9w34x+XsMd2OdFsYxQFTALDJwatU9yvNQF4
ETmoDUSfjoshhQTHT7H815j/Bupak48ZctiA19MBlC9u5iveU4bM6b8FB3YLAFB4muuBOFqb2KYI
CygeIn128rkp/QYxlQamqQdKaXyKdK2+UXazrGtMBUQ+twBHuC3kLrjvQ3r6D3fS0TSf2bDkb85J
lAOI881owNpZYpvTezf0Tgz4FhNAZFOz4JlKwNOp/sImokLx9e49i77rlYp5wdGxa3D9xjtfNTD5
J9f607bdo+CfVwUzKNDZgG38zpOp1opA5Odw64/7mh9PiCY1N0vEMBq7AN32gDEVWgW7nhAa0a3p
MD7w+o91VkBvyf/Iw2sbAnryYMm+MIodfSoeUPj8d9grqWoiL/P6LVmjKEZSnvx6b1OXIFTTRWPF
SD/Htu2ti2amaQJrZCMy3WgTXReD6FgxHZkCTpYQEf9s4TnsLh71ui9kOj7ybjI/ADXGR4VlNWLY
7thjyjHXXyrycWueBsqEDYJyTa3KWv5G02SQfjG/xSXiLnBduAN1ZPmLoWk3WH6Hl/ouLY5iimhQ
hW5lgT0H0WnUE6qgNW3/0W0XERU0QBuru2qollIflwur68FgN1zHiChMt2BLlwrZAgzWWC2XacDd
akKmDW59q7iuPqGU1YPivUGmcliiiS4CYkYSee0kEDwXODPCKJN6A/sPWgG0gS2H3yu2IHpGBV6k
gxMYXIQGaXyOq3sYikvZxEdCpA//Dgo5mTixiY/7JkC/eY8i+uPluZ52l5jc8VZZ5UtLSDqrWyVs
Lo2rBhxyJaN6444jw01Bw8jCElJKXeQ2V5+1A96nCutXIRJBKAIcixlOH1pipvUWHGnNO8sjj0bU
ZiNHMqaq6Q/oTvuyS1+4CiE8V4uhA4L8olXZZakARI2eSSN+J383FjCC/ntvWUswUG65iS9OZV9L
oOeE6ilXl1nUO2EGyuoCIRENsliiZ4Rybx08GoAmIM7DLnc4wAIRgb207nkJevbdNGSl/LS+n2th
MTNvCUPkjYXBjcUGkxl+xSuuwCHJo3VI8JRLHEkWP2zf5VcnVvho/jTsUsLeh3IvLRoiNODLv/VB
TASKAhAwXdKCyHSp3x5cweqol/vFxzA4SgTGFLseM4n6juNpB5qrV6WhR0pV0/LI9Ktxuf6akEKj
27FJhCaluNjltnHngZSPKb19HOFvVsgN7F7ODcVbWMlyRo0zGMSoj0qWYX01Dxyh4y8578vQYmpM
fVcTqt/xnyv6Gq5LvbCfMUh5M3RFUkEEZR+OWsEFdtw5CRT+xqSau4/2kokYo8h38YNXysSPcdvu
iw7x8i9xTgnU4gCtsuZuJtbdMlWor7hMbxk1gUlE64zXqDlefgy9KN/3eWE5hFVTDZv45PUIEQb1
SEq5gNRejrQEQaPu5UALGrzhdcBQUd293TZUtBpXa8+I7hm9/9tX8Ks2jCUb43OWXsmI9k0yo3jA
LrBY6hfz4qwjs8kUSoVo8Vvet68zUZxgP60l/yX00MWaylwYnALLCjScHcgmXIvy/LF4nciCL44p
mhZzb1Zet0amxlTM17RYfQCQCra19nE1+O+VPDtFWRdxOG1TQwCQj2UexelyInXLjGzodB4dQXvf
ndB4VFxR5251Y0eNX+xysTomiCDFsxB93K/h5V07AfM0+42C6Kbz1j8OuyqK2+3B+OniuIPdLG1S
+lqtcw3airlOvSurUFa9/LeScY12sgG8WdWCyuK3bcoPrY0i4RKRjSzfoOZaWqicOPyuFMhdLypX
SANBQPV8+6GkEjUybqvK7S8d4xKDnE28VCc2i2HDL711xqDyzD7pCYeIZYeKAcDxWWscsazX3KK+
EZtxGpETRR9cxrhOkD8BQbg5YAowWb4RZo+Pp+JR/DsZF++Bq6hcILxB6Uc41Nidwxh1JRPD1UfG
oBso21yCeLFAwvAZjlDZvVjGeivvYOFJ5x7/RyNg6WsfKQ+YPXWR/BFwIMsBAzzNu+UinxIROuzf
752Adk9IfcLcAMtCTzhfO9uhg90oaiUlxB/4LcWEIN5D7n/rs+Qci2rTkG+yG/pvWeYj+nHckSZZ
dYN/krgLutY9vZBUv07OhzrAaEye0DIH2teN46vBelfStf73qy84qGSpaqu0MrN0+tzryUhJz8RS
ZDbedYSgfFL9axzVQ7NW9Dg6Z9cgd0jih9YSIUoWip/zvX/0UdqmCVu4eOadSUCHMNwmluxMSpvq
QipL4/z1wt/XJhjsuDKdxV4AI2X+kmPuBcYVbfwXvGH7r2XJqr50FpfnvvEO33qqG1mOhPM5vG9f
VqsjugxF2MU2PbY4tMPwUYKmZ4uC9QhPJjBedQdVhWDC+MX/MOLyClqMz5GsOcdp7sS3V12X2R9S
SaTFfOnXljlSkwau2WggPqNbN+Xnd57r+MYoc01qSahHVnIj++z9w/bQGHZHzeCJ5K0BiQfE6/Uw
xEEqydc7Yf8rt1F2e5os45bL3y7073NCs21C02OynfWP0NiaAWl8PLO19sbYkUXTDuNDZZNZv+rd
g9W4AP5fuZQWtkIUJlejmxsEimXrAKBA74w4nqJcIMAsDsB8uiygq5MzTAyacehKgAjImyEhEcmA
Zxq/ADgbnBGwaXLWbxo5QOZ7cfmJFH8i9a9cxToZ9I5D6FsworzSuuyHL6FSVJ+rjmQjmUD59N+1
p4KIdiVGR2b/I1phkPgue+M1wlvRcit7eBlZEWOqX/2M/h7Up80k3O+oDP3rsstKz+Qsi0VJ6jNg
qRfhhK0wcLGNNDgzsW1Oe0InGWKlhbxPniSiMIbd956nr3JBWM1vKOPxUEN1NWcBjJX4rHe5qKNf
VfYdOfzwqVDzttfRIUgtA+5gqwpTQGMDKSC/78OYY5w0FuxbhKYtcWl65fpn2plRsiv26IE3numN
l24jv9f8v47H9dsDyffEPBdQ1jjZ7XU525nQA9i+piudXNYhU2hb9eQaje8jlL2gYDZpFZhoSdn3
hzskh7RzAi03d02YGPFaNE+u5EkOTioYfF5C0581l5gMiP9HBVIj8AYH6o4WfuipDXDIPfMR3hXm
elvDRjQYsNAdnKu4PV5az5kzQiUPVOr+rftjEnwlR8KdhxinBGVrOQ3jd2qJfGm2rfIBAYwPKq+V
yEl6kjRH6zE4WOEMyRCXXfilcvXymBDYdWiRBwTGK0bLizN5rJuWwB0GtNegrDY1TXobj6db6ri5
FAH4Ku0yh48pHjEs154hezc0O6sbagQdwotYLxIbPyhvPhq8d5WiyhlWFBDEFktLjlnXAEcpJqCC
P44P/RHoRa77JAny70SqCdPPD8873/12DPzsQ6YZclF9UFQTJeL1k2HwuvgtMFwDa3btjMLxNCAa
zBrZhYHWpgCMpfoC6h8eo7lTJ3ouxSK/58/s7I5JPTJdk6N0CfxV01pqAprpvoEd/IFyUYcIMghW
ItmnyBxmdiXRsiyKmKpYwuFdeSb02HtbUHCfTGuwHBMv/HAVT21+g4M2puSWBv6S4to8fOPSZO9z
rtYTVFSBYD5lyQZpFCN048vSwKpRRXXWtPrlg9Ow1lqRCfLeMTUb9iCq1zb8I2GYDsPL/czzs4i+
i6DnVDq+rC10Bnb1fPdrfy7aNqdjt4N2zHQPJ0Yz/JINXXbHBAD3FN+wZzUoIXBl8VxoXDxmj8Uw
sUDqwuXVltN03TyUIpaOsKSqd1LZxcD7Ux+AXu5PHEMOMdg7C6RzS+8TsYRxMdgSX8eQUGvGkPCH
s09siLQdw7s0VYJxGuxTsDmESw5i2DEWYstue5pU96dsVGSQ3/0neF3J6utno3v1Mx1zvQ/pRJuN
uuJjtzFFEBf1uHY2aCoMiwF49jt80JZPTKbJ5iOGkXu2sovrQdVu+Z9Et0mty7mxCZAe2YBU0sWP
ycToDXd7YFdfvmXO3vMQFm0wYGPpTAXLKmrSaqDpnrS95HpnYzjjS7LOBdsakH3DgMcOODBlAUlN
z4mmLadqqpjVnIrUeN5gTcWhOiDiNZD5Jy9GJoTVzqNt5lxE/8NT34HSdrMETLEk6kne6dt1dDVt
y7egQQUFc4PyJrKwVIK4JcZ1Aj4qGzwAaZcUFQPUCgsmF4vpTJ0oiGb7JbhNlV7MTWBkTAv2wnwD
WtvkiiKgBe9zXDKFS97WxDa807ZoaTwnvFaX6VcdeCtn82I5o60CwFWDYAjJU5hajVQ/triYO1zq
obblWv3ZDbILHJec1aiYXsdhPWaujO74FN/S//eWFIM1hBAS1lVFqxpvbSUat+3ArwEL3nVugPai
o4V9aU2O2pwm1mc12o5rYkmwCPmznLIVQIUZGVo4M/iTzppBq3IZfDq6xt7YxrgMN/MdHjvOr4UA
rzeDB0L06YQAGouwMvKhEXXO3QhaGwKbaED+/PMgkpKCvqNjDYSKikKlf5LUK1JrX2PUOdhi5mCN
m98IMKjUfyLfvMd4XaQEJyE78HkxIPB1GzgNNgsWXi2s2d/gYunEzOZ0CUSVGpzoF3n3+FBSVYR4
dl+eT5a7wP1a6Bizvc6aJLOCUKSiG8Rk+VCWwmX+GDdu6/XJtS+FCd4fdOOuHqmgbC0GunrLzJyo
IaG8gIv2MC6KYOFWh8MFX/Hq8ar9TwELuIuqKprbwr9S1qKew/3INH88Ka6dmrmuavfBCzmeddlF
x2TjVPR4A1Tq6eIPTs87dMpMM/4gnpMr8l8OSIHNIKh2EwQTBTQXAlE3yWCExjqJyNQS3erxRbx1
nIol/ViYBWH0z1ni1xFgTHRzwsQ4PvK7ihyB3yfJpshIWkHYGguzk9uJEAiGEZB0+QWANtvr4cem
dM4IRLMwED8ssFKlzu1vRkhXD+JLflYLy41+Q4riJ5x7CU9M0nQuAH39tBySR8cMD8hAqRRE3rnW
U+rJ3bQO0BQabK1OWj/7ql1o7OmbdBTgeUNdPB+Me5ejgOKkfR2BxLCPJf6GzR28aktKMY4E5K5o
3M3JQ9kC7AdrpORnKvnZ8O4tekCIwl15ot3bolrgM6hhIJVD0O6goZS+s2X/GIgwvxep1UErPJxP
yIwx5MUfCB1dcKCuTlA5wUR3GPxWJotJMWDegX4Ay8Ey9Y9xtWsjWLEEgSuDe4tmtxSIsO8MQ1EN
xVMmHEaOqW1LsWAeMWiWfwGjQuSs9lDx23sWFExnoji9Was13aqtUgs7E2x6d9hIeS/7/t5RWbVn
Dnj4YXhPYhWpesKRvehCh+4TD8+kaSbOsy6AjMIdnCyJhIAGIQHlHS7w8Feg+/nlU7jBtd0sOG6s
frxRW5Gy2qHwo7o4ICi/lkPGtAmFyjLsG4HFqeNQi0PJvqpBVaO6W30TNlIuvu8w6WmE1WH/5trD
zJDAncSIABXc2tg3B0899eu7LVEub0tkpahSuPpDVXS3CZDV5miY8MnL2KSkaazWCEfb1PkJnTgl
chuXJLPnRjZWvgqDA63Q1vd1v+0PEgM38oOqTYB81kPo5XagBflm10nqMjef0FVN3JBKg6diXqLD
iWTCZSdfXlekxYtAVTsjlLqv3gozgXBwAnAp84nN0LFwObLZF/R+MXOZ3XOJ4Fn2Oe15/VvObk+S
ZJWJdyuW/ZSV0rcPl3629hFtfM6jtpKSKca1zAR8EhDjD4Ucf2K2oK8XJnhuCYKTwtijR+4xm6AK
FrADgEch1R7nRaXWsnOtkHPPhptOWPf45m1BSHkqpO05BzmnNSW4tBbwQHGG2LfPTZrseSaC8wN/
WmVxp1V8OzAGSWB47D4QoIKOBnGWyIJu95B7q8dlxupN9mQhx0QR6zh70a1LWcJrLnJ1ntAegtiS
brVSeE+kDkPYsaRUy4UVlI9THvgT2jCGp4w9U1QDZ7AJq0XOTuPdUYcptDwBBAMGuuah+w4WrcXY
am38bEgQeepsHqQWkX2c2e/Z8zE16MZQrQOhe4Vop7RG9uGbzOIYHPSTsx4kXEqs9cwmExdzDYZC
21QbJ4dhXr3pmyAZ+tf/ltl87KeXFuBaeQepw8XfXNh9kWQUROKdm+LJcbyXZW8ZGcDnCGq4myxO
dNpi4uLs/lN4RrWP27/nmWVqYIDPuC0xpSOURBQUxEyd9n/mxdukdiIbBkRga05mUF/3tA1Hj0z+
3LThei9uPU2yTJJ6HBczOGBDjf+R3WQGutee20fahb8gB6bn4JOmmiQ927Ngk9gwhLoo6ZyjGJw9
2aav12/QFJe+ZNqZZGPZCMNmSAG+sTV8wIKEp/DhzyAtK8z8IE2zVxXehICzVg2jIT48j358zCVv
OUXeODPUqWE5DQbR9Pt7nZjjoUxmuPhkogZdPs3YVvcBQx1UhUrgs0ZKVL9CTBINcpidalbIlbJG
7+cLG4jc4oQseOIAC2iQDbegYP6Oj5iANig6EjJE+pbglZ9un6NCbkCUdOxmqovoLPN57NoBPIlM
f4FMbrT3PWiGW0Pa8E92lIdcrt5ldLY2hrx2v8ERyALgp5IhanfMiXLw+MWVipcG3DPQqppeyx+H
LQ7ybf8LCMp4XtO4sHpP68Zt9ubsFlmnOFKV+cTmBZmdbXw1IB5VXPWXTIfJ5eDDaqXMc6GUlqXE
QfL3pFl3bNGks/1O5SCro4qNqWabn/4Qg3vM//zfQdyV8mfGp97XXfA1CZofspEHFjZHW1zXmUGL
kh5R4VhO78GeWxZ+F/NUFd/nk8Ucr7TJNIAVHBUrXVYvTD7syB1KyWny8BR0HZdLDNg6mvxoLI7X
uUGbt+ti/IgrEHDcjHstjX/Jj/oMfcj3hcI2cQ8oPyTUzr1XJ/PZKST58W6KKEOKqeqxSfz4maFi
jJqCBUwdbnI4qNe2+tek7C+6tK+tFWY7UB5oS6TUtI1wg0kytwWAxRTK28hb7GOb40sfRWsLs3Iy
R7Fo/Ehm64+JL78XDuEmSVAU5jwlE7pFALbemP0heaLjvarNx29TQ4hm/iQZksaU1fgzJKK9kD4W
cyhP4dlguhHzE+R1SzsbJbIhUgmRB+qmxZ2mYzj7150S4lb4VxbEF5/Yq8zY3piBd8qHvYNP/mNY
Ezc3qCcenOTntaO6J5eySPcZN9zTc49J1mTlYVkbIFc8bDMbN0m2+MZijEre0IWe6KePCsHZG82v
fJc7KOfv00sU+HgFPNWdhNVWfAC/zhP5YeydJlujZgloZerOrfeb8Icl5l3ch6fOS4U/5p/mXkyN
iJUAxtl7AR1gdxSPxm6W+MF6q8gEH762d4B4eXSTQxJHoTBjpMpFJJqmDt4CLMVBjZMzqX7dTIiX
0oGK3BblanctPqr4tmJzVaXshcVtfx/nlzowZQollmxQhbJysYLUdIoBZ8qeIP5TFKpsIjijsBbm
xPRLpnYFfOAab7nkPIgBGUI33imiCU9/3uSkqWhcRVRHJw5cIjpaVZeQWVnvWqh8iGimqbt73wwT
v6iZoHWWxEbxB+g2glo6NMnI7tynSG9cikPeJPA/ilFpJ7cqtAZ/9gKQppMPMocv7f7CBTMTIc0L
i2uq+P6yUnhUKLB/fECaaJ5tb3p68VBt/1iQqUbQuQJOWLqwaTqIKqqQw5J1L1G4hrt0KWKs77Gi
7OkSsvhjwMUzhC3anffnN0zefHTEkSO1gDS9/f1c+FIoHhUyXO5fvKeRpmE6Sj15HoDUi4rYzmuQ
+WPEhoksXhokAlMecf4UOo5umMrfoqdTq3FiemOKOM0xI/VERcv6cwVk6sxizlC+WwqmM9Hzh13Z
hcWSzBKl51z/pl3TQs8WaHol79e4r2Wk5LJHKs66ao4NTf6zfp3PwkbpoXL9K21rFDhh+zO25BtF
h0NUU4j/w41HLo4CfkTWNtp0vtARXdQeVDnvMlW+9evOchkeJrY7BNUkpWtuShw7drWmIaRpybhd
4xnUtHKLKR9FYly6UxWNPsFXG2IvklTXRbWIbQM8UveOzbhz23/3PsMnXrw4+M3eTJFw0XH8t1rq
bfAWWWanPKPrmrcbfXuZsEzI5wJCStVM39Hoi/epW6fjfR6Vua4UlXjfyYm43noF/aaETGc1e8Lc
RaK8hwcUtrw3Vbkpal6+kNwGmHeYTnU0hMD3ovugLQuv9lzas/+EM8Vdt2nY1oWxMw3NIKA/o0OW
lPU/UNiL3pqSg+Iknvbn2CKBOG/RQr2S5LJBcbTHI49qJSVmEd+8bgy6u6TBD0vvaYh0gBwXAi2k
GmuOWII8St2+JgCA+zTJUAqYRaJllf2viKabeaXIY+nernlCDIeRPoMmzWEOwIfe7l8u22AyqHZo
H6rtAx9GBBaXlL34LSgEHNvUVvQRh+NPU93ljar5Wp0Hg4rSQCowKvJsRHFKnPyr5R2yNDoPylWe
zjrxfBxlk2ujVd2FGUS847ULFV6XMv27Vcd12i7WLb/T2AxsQ+XtbZwTbbd4pm4Q4efPfKP53kvv
lXge1zWPLzkvcSvMt8bnz+yo9VtKjavAJ/NY1SMKydY5o7ZeTb9rcc06C2/nL3ziZfKvtOFQgeU0
yICPciQ2bDxO9vUOhYqsJHzgoXNPbj4OkUwMSbrAfT2z+dABT9SKys1UAQ72NTZJq0lWaY+E2WB8
rq6XZTevQdiKwZ8vuRaKxDxXU47cU91MGZxqWVYAJ9O9vwvqJwHlIAfPpjxeR2POGFPHIN7O9bbd
kGAXg87zHeHGZ+t7qn1gy38mS38sEjAItHcqqUTy6JFm29kd5YzHNkeX0LjqnoeGR7YdeA5dH6C8
KiTMPadWeqWCAAwwP6PU4pEjiycXAnEJcDsDPkRThMKDkofP5S2nM6sITN9QGNACLZDSntWX/qJm
+Tl6PXU+rxFs0iG56zDg/dq2UOG/nq0GjCv4W/sW1yGOzwzXWUrbJYtTPlxOkxfD8KTgHWQZHmHv
/p2Eg1B31y39kn1vdx4DI/VlxfNOdaDfJc0xHKnws/tGrIkTGAIjyoLwhIHSMX7+5Q7TzrVvf8Hk
aV44hZOTSsmll2S3fjE4UIQkjcztJLWMGNSXMaia4EuZyU+krn6RmC2U/ddSTyTSaE4koTaFJKt5
pROpRAWLtVgvSlg0aqzGMW0R/RT1RrKrNn6MnKrurCUoQAy4Tii/jqcWoAnnrVGICvUhQMhIQe8E
0uyXc1e4jDA567SKB98a6/Pjd5nn8HuvH1UZESutL6k6bx/OC78LsXJXLJnj7vFaYQM+aKeRFATa
9kqva+rMTP14WzepO6URPEZxwuTZ2BCaH61ncVHqKVkU2/NisJ/1B1SgcK5+9VxVx4M6b0MdjV5O
grK0pRcCWx2xGGu1wFs+R3IYBo/Nx7vjliYycsZW40vqSF4xquCXq2hovjcxtobSD//S/GLZ/5Bg
jcxSLtfAGFqYkheAohH3OMAFzg6ekGadEvOKPwgo9mI6E6xMeC/lb3XrDjcn6j6ztr9/Zp058zcL
2Lyp7+2DYzTWqA9VVaur1D5PcSc62DOtg+C/aYq2VDTEJQl2+MgYQaAxmYQdexHhZjwXbF8eXtfN
oADHPE5Bh3qns05ZiCLB8yyG1Z1V8hZmj4bOaYCQ+qAX9bUIFpyc7wyldMX+cIaQdGgRn9iDVWhr
Wv3fERDFzqn6V7jlXJByA70dlqd/xzk0Nn8mRYojGfj9VCrcflWpqAK7DEatS8NMdDRG2fSvMPnG
ubkiBug3XiOKKVGh8KkRw3mVrSO+56e7ecWjor9SI26DQc6ZOFe4/ZGH1hhiItNzMr4XWfZQZulD
qG82usWAN5oiT5G+qIVqq01tcu3PPyOgYFm9gxdjdAKGUIcmsrTJS8O6HUnGj756beVxzLZn5HIq
4nm+KoCsFZ1Tf0rat0PAxmZeIG3fODZEwGVs0q2RloGgyZOMXnbekajm9jwbnQGDTEz2DDZHD+gD
djhz5lwEGxbRXWlMnVmeNeAOigjjDcx4MaKDNOzcF9g4lpd1bCuU9sSS9jFxG+DGveU6Zlekokc2
ZyWk/qCUYnvDyI5zr/KUgpimck9shIpk46+qzyOBtTDXTEu/ZgTzKEQM26YNh45tg9afO+ywnQu4
YbdNgHWddpYCAy58o/g8fliUcWMIwJgJ70aLGtOlQMSKhnKfw0JTGKcjIt8zGd0oprvyp2rLmQZS
UNing+KYg/jqq0QVrEW58N/64WHQbIlEfyHk8UX0REjPi6I90VG1adHWcEhApnvdAShsS6/vqryf
iz8d0UPUEWUymCV4gPP1M2qK3rt912jwOnR7pvkoKztiluNcKz5iAuJuGk3ckclzb2KqcMY0L5CZ
QQOkG8r/tMptwsyRpOW7xLbhX35TO/8WOASn/6HSRBkjiwjX2DAkA0MwN/SqLs/FJavmZptuRmFT
cs7Jk5wivhPCbRGrTEeltjeSaV1909abU08xSUlHa9LVpCDFX7GoqbwlWBUMCFyKmdY7tLqok84J
wManIWRPh4JLa3/e47ltMwPAbQ5MTGLHKRZ5JrTmPysnK3Q3l+gS7zXL0CQyisJFRGiDt4FGkXqb
emX6qUl0U2MZVDi2RMNjfPX4MtTDdSY6+g2D95KamQk5FySu8H1zyxgliHHTv2UqWVJ4mG7w26fn
kXG0ActEuQpMHEqQ+/CkT9oVucFS4AduoJHt230A9Ehr54F45rqPfMZMGgqiuAESNJSf2zxCspgc
xDtTaJR/PqfViO+SlKv6UqF6H9ZUtnG9T7buBmVmlRZOEPStyNN67J41nadHLsKVin05vZaEtRMb
tmrK6FSnumsj85dcH7r5/GnqWhayr/p0LvMHWHuwm0PcaFIh87AqGZf27VQ+c7PVLXdgR8E7xwO5
vZuNL6U1B12zcrZUZphTxStgX55j7jFFSqEbavltZ5LKDv+FKl15iIzfUQP9FfOgUzz18Tr8Saan
jJRqvAuA0EqTeHxVHsmGimWn2XObKrsbLqw/F24FqDaV/HcxXJLKXrvUv096HlADopM28SIYy+xl
p4gYp9Xh4ZvQeyYpCJPISP3P+svgSN7A/E+XU71sIw1WUAf2IKfAdMRwV5TAhhw25qg5sGyZ8LH8
NX6cHbzEaHO3cQo4CFopv6S69Gt/MLubH3knKacEMmpFo4oeVq9CwysdN1mbrBapgAH/Qukdghtw
/Kdgpl3nvOKk25f8XgWcitzhwN0OvRS3s49BF8JmbqYJSYkNiRkMHl5yYQvzrLnOiW6RkHpluJVi
kLPhpNJYkYnwF2iRRb6Cj83PxL1SESOG/ONMvmAUtv76sax0C7tuWpizVRMAWN7Gml5QuAxso9LH
uR1VcA5NFWoXNu0zSi4Gw2kAbdSmwcP6GGl7+tYCIWNswyqIZ1Doe1l6xdTgdwqAOYaUAMLE3HVa
9AFK46KL6xHy5vnK0g0tU6F9GUOSyXbxL42ry17yVU3DIxB82+N8lAk85SpbY/pT8HXPkUm6xo8o
cYe2Eu9XXy1DOI05JGcrBoRpF1PlhXefC9YH710u62FZV6cgCROYT+z8Mym5ydw8CYW2UTX7691c
jYbVtQ7FN9BletpJH1qGEtKF0ddXFX/3tZGvl+uH8lhG5B8TshBYoS6smrD13AHbAp2MN4OCQJ8U
WQ+b3bUV2Xejk6WO7iq23wnG8pIspXj8ugZNpoXjwSVfKHMjP4wVYHRzoXD3znsHaiq32KiE2tj6
o9tz/OMZqp8UkYrrtE4nzwOTm6VQpKV9jdCHwHuZXsH/r0Iz1pXAa1w2/HtYKZuUct1kZYOo9PWJ
qDS5Rh0J9Kc1Sx6dO+fyJ1ElRq9RH3fEZT25BLX2lpUXPF9yQTbAXfY/AZDACeGQ6aGDVHCyZAuE
A8eI2f5V3EzgYJ1z1nkPVXP4MQKC2RMGE4lVHTi28xioIxFt2LPP9quPXEvzVY1llr5UervZIGuw
Q954VCPWyhUbtdc0pu5NESp2JQzxNXP9EDn0YvDl+gZAH0xecS/MouSp9u0/OOUIjtY1KF/bRtU/
dViIwPlQ0mUm4f6O0m0yYoVvr6jHmw/kqfXTAEOUQGFox0IOdPdw3vo715XDoDalR0EmGgLeEGMz
iN/XFjyZN4g5Yj72chklxOKW2fsq6ExAITTU811AISF5m8vOvdNgEDD/2HdCmCNkyGZ42yT/+AW+
b+f6J9bRv/Fh7nzV+lWywKmJxN8IoejtAPWlJVmq4P5GZGtlTiFj0Yfk96PTmVOlbODxAxWQLUbH
3WrPfZoE1q3wmk77twmF72fb9H0Xa2LbXBnQ2ZIXWaAghY+buTxVRP2kAvLRb1NQcBEnU5CgqUHF
QPPfHTpCCzPVlp3XJWpXNCoq3URCt/XhivnbnBVsI4G56rL58/ICDJ3/d8C28bcIZFM4mbxgtmfx
x5XjuxpcL1/iEUzSSDiIL2+RwitNBndCILqzJx82ZxD9YOrjxm6voat971577PU9d9dcpS+iiMcI
qIdwpDIU65aOnwqJ2tidRQQpESJ73d/W7+Ayf5UPbE7OuLskhtKRoIlxul09PBkn4W7xc+BnTTNS
+nO4OPD6/r/s5NURWjWNoMh4pA1INcoRNteobKy5ESQlM5UsAwZK3yLisnCMTfAsbtgT+7kSEEHc
JLvOJANxxB92ie7qaMUxv2Porqy6VoFFarcq52N16AOJAcd6+nzysTebCIIRYMeCn1v7Z+/gskIm
u/zFRwukpy8w2ScFYl5PtXoFGjY7ipJkFLOyTSBsBsGpyKWvqgcpr1epErRA23RW4Xts++N97o7f
rgcgOty9n9tjpykJDu3KADRFufQHgKdb/GbNqtfNWSJslWqdjy5kpHs4QVm/2nkWEfqBX/kkGTTY
053Fmz2aFk2aZeBGdD/960ZLhmlu2Go8w6qJepvSQFsb3IHQ+ni3dX6obI8D+iu/MpxMl+HUZS1y
5kVprMypS1oL2po2DX8GTBex77mtw/tRRp/Yr559FSyUrlIldWmU5T26vCAJvodQ1Tw4LwiEiBP3
pOubgG1GNYxvHtuJ2wzNHtYUDmInNB9kwUrEDH3SmL0bGosOGP/eaBn438wmNYehJbIO0vFPLMOM
huSMAtwra2oBd3pV//dCut2DLS/jcaL5ry/wL/RrDd0XUYE0xndAYT36mj1wFytSFJH165VzJkrB
HR1nPyuNVaYHQ2Y+TPNIw4ai2MxiV0/uZQeMuOgNBot/+Jcmu/XW7AN7DnBb3Au8FqUDN/58BzZT
klpZVfEMXF0Pp+nfNFgwBH65Pepe/VNm5Jbh/i2yJ+5FG387Hx/dgXKXhoI7qrKmgUhQKkUuOZl6
sVxpTH5SHW2vM4yipOIO5RF0r98VQNJbjF5PedjcTNCFzefWsaAytft59dk+tYrnV8RsotI4VxX4
x3fjnOm4Uid9XIHUhY+Rpd8COXxdMewMhERRn49VsTzqa8aeD/vdVe6DtMJqXS5Vc4/XrX3vOzkP
OKBKxBveQRPv4qgs9phP5EpIQqhiBy3tjznkbPHf4zvdT1LvC3/iiPpM6Gogyag3M6nUc0WmN2UV
Mi6Yty3a3vitux0IeNRYR51Q/GPKgMgjBkzXi8cu9LgandOhHJ2tkw6B4W/jVVuP4KcBo+jcc0ev
lrw0HPL3lYPN83iIrVqCVA8mqmel/3jb4tIVZH/6aeepIhPeLH1QgPrJ2jGfJoTNvmpBOfFWpbE2
tH/yTfmN4Ie6X7vymfOrG/5GIOcymMRqsEalTq/vpBrSLfOUebYdqPUuxLOi62jqnocxcC6CDo4I
8SYprs8yhecPqHr3+YX4UbSuQt+jP1bbbjb5gsg7xcB+3UaKIAuXnrNykg5lrpj97na704wkHBG4
+rr+m119skdnuhnUx6CFL04aLFvSPNvrY5BJtmadkSE/UZA+9ywxk18+9sDYdKouTtUU5Lrq8DVM
9kzSZXZe0Eis0TzWYndgCm0q9tiKn2CFT1BUxVwnF8PTrK99+pkLKbDvjltdhhXm6EmsDePzFHVL
d0y8YGbyytaIkjttD3wsn/1j/PAZD2DPJX/LJVaGS9YbeyNfTgp9gAupLT0yZbiLpQxd0sc6cMuU
UjMhSdlN2IFwbLk2Dbiqa6vQgYXsXJ1vTETdEQbkkymgg6mTlrUQMghWhuvwaLDni36oe2WBS6Ek
MREx4JsR3dPEeaRh/LSUAgWw6hU5X9wy97vM4kN2lfEr7Blitp+Fug5jaazVfldBuVIdEZMetxQo
OqZaPSsaZrx0rDZ0gKANzoWibnjNa8KFEfpXvWu1LzOFtnXCODOwBqsffukIAdqw/6uygF0rctMW
Pd6RySPnYEY85flz2aitJ0CCH3Co8L3I4tlPR/VZFTuCqRETZ0MvK4hT3VFEKZUoARKiGSK4b7kW
w+UZT8XVFwu9KsHSamHz1UVO8RkmN+bURxqwgOExlzCTrvwnDT5VEYI/MttSZ7GMXuHk0EWOX7GF
swaODHqliDtUcb/7VF5+xsZRohOu0uSUwDQS6ztxfs0qErZfkpOD1xSfmJsKbFnIXjc33Ve6j1QW
4FuP5FWjPN/VTjhJWVEGwiadc7CDor7wifWYA6BbOG0cJnYWEEdLtpbyac7RhCXaAtjO99iNuNQL
z/gpPvhD8aso5gEClbRiqm66eQc/Sb6PgS8KV6NEi6ZlNK6Emp9PMXIVK19Pqvw62POupUOx6cbK
qTYzsrsibR+1yQuEWAkVLgQcIPkQAGDUkOJPe9nOAfTlW212ChBs9911q8b5BBYeMttG+djh/uPh
LXqmiD9N7uvRf9Tv/eymih3jY9I1cd0BSQuh1QNXbzvr30i4mDikkut21i+PmPc4sXle/qUTiI96
m4Xu1olf8qO+FSaSVD1ni7KjYZT241S0nzD9VAY31/ORA4Yvh/bHEZgbO4tRaCBiq08RhwTzOKbD
sotUrsPYThoT7pMdNvcH2sVZWjlByU8kpa0DpikqBjnW/5141rLOe4ylLsnFkqKpEImhpoqTqdfP
yl0OlROG1kzEDkbEZ/DhN3BSI2bBM60X4p/3vh9cdfiyS8ckWBBeIXbGwBdNy0TBetJU+hSKwm9z
R3LEwvaBiE7Ty5ip37kv7bfEs+6g+COikOmvuclgGRBIVyqFP38PCUYkqBXDuviEXdWjEZcsovgR
PIiP1XTHYbbQrkhoJxPxr3org09l7cHYm7aSDQH6uFrooSmBihWrfb7TXLKckhGfIE4gbUlqhplR
uscX1RCpstpsQx6sozXVr/jTtHPxDpzTP8/pCanpPIFs8pVkBtEkhQOGlOieUX/xxyxC7rce04oO
z4RnhuRP4PkNN9QolqpdwNwU4kEV8t/mMpLM7f06kM43kU4fEdiJbdzvhgNB+71895xRqJdYy6Xv
kji/zdccmhoxs1JzWy/PuczB4EFrJXBYbDrO0aj4CW2hJr5jRDxWojCSGEg0sDAhvd9cSUFLdZtv
Q9On6p8PmtMuknwThCqAMZCyPJudSeiMVmYPN8oTUZjBJX/cjtERGxrfz1OhmiTjx0zUcCmUzftT
5p99Mufnkv0dVsy6SdmB8D5QJLUnSFaF4rSEN+SFio4WkL7CJGR1m931p6IIxetY8yo9LxkJmSRx
oI8myoPU40pY+MweC1USPkJuOWzZRmnu0Rj/dR4ddl7yD1cJiIfsoZqlUJLFI0rtVbsbVCoqXQpd
ORcKwwNofRWTFgREtbcEcdTu9TUSJCkiCCBu9c0YUqFxAvYuBEvn/qElUoSgqkF2r0TgfUitQCr9
2P4klBOV3Ilet2V1yNcvG/uUdFVpI2zkC7MSLtUeAjZYtyf+Tr9He/LFkS4A8B4Ne0skB1E1v8pK
k+8R9f5fT51DiYmLrB7tAsGMaoegEgKxfBNm1BEv6w0ZjzCfIvYs5f8zOo14e80FLPY8cnJ/V0aD
ywKEB9Wy79MgUcYTJMoigaOKv0F5yTgRAnvK9OYI8E68axM5jXJtzlqFtYHfFzyDsS2qKns7tfm1
tpR0BrhQvPTfQMITGKisGUC+6wQDYKni86zX1yX+XzqeL/BENnwmisxNi1fLqeJ3LR17v5nKA8wa
ZgtWp6uXoGWX/lyD7EpNcqvqWXd5lr4DHaYuuu3xmY50ZTEhHCUgbb+EN7rvVk+zZGQTHtai51gB
dtuVeaEMozYtWXrY96WbfjtqkfG7LXUXF5DYxpqV427L3nm2EraIWjZ/7WfKwjRUVwKHpEuDjH9x
k5qsBXMdiXODntZhs7JVv8NgkCgoqMkM0wCold1z09FFjfKgW8mffx8h91/8+vSS/yldQOGmoBBc
itk2wwp1/0GtXBeWBT0CCDyFPh6kxN+yWZUNhqKB/AgVtXG5Xymo6ckKXcvfpFAjfJINguyBw0b1
7nbhROBgguaflVyyquJw/itiOqz+jfAHkNwv7TvcE7GP49iacv6oPZgDVHDGUG34P3n8Qd9woDS0
toIO6ZVj13aYuROrmRk55yPxgh78ilon+gMPTCSpp0evf4ktH+2hBH2cpfx/HwtpPtTLvyDVnGUX
icPCQ5BpNHkEtxv8eGUz9RmuYImn22RKrb/E9JqQNV5oPDurwBWtmrCcrXgJdwsDco8nsEmydTzj
WXZlLb3okmXCpqNNgQrZ4azzLnRJ/mk7joHMJ0TLX2lGco+zDhShYQH2TRS7h+1gf0wpb0iFf5Ln
xmoj7voJnBSwmemN3HkGTPJ199CpduD1fvhj5LLzHkM1kui1W26YYQUSdlzU7RaCyXiGMJWEmrK2
rZS3Phc193auIbg/yxSTU72eZiJHUVC4CatD+sicnXoshgCSBFEkCVyJOHhNltQSal8LHzoIBVdB
zHHWh3InHV/do7/quBGKhrpeRxkDGq/6PKYbMNs7P16sxlSEwlSYPyLBfnKfMpYl0VS/5f0PT6D+
+miFJ0p170DEBaGOGM693eshYasxA9EejeQpYxjM7gu1PLThsI87tsM+Pb7FpgBpfL6Uh2Lvx7dd
ooJuzdHvEsK56Sy0rRjzX/+bJp/FD5jlO08iRd4vCaIWlmyOMUmA2qPML+0JCrWVyLe8OWem8mOL
qls5IEpBix0X0jY8iPsTAZhs5vNFEbChRN2xwNAepfNmBrMoQCkyAFru/vGy9i6VhbruO1T3x3Ck
SX1m3DFlccdrA1005NfxpoBD5StPqTNkfFGFEGKJxZnB3pp5HpsPcH1saBV4YXhfk99hmPRr9ie/
ihcHARN13lg+FUItiLvV4+Cykl9fUVj7Zu5Lx9pDRP0VqqwTgVbq5kC49ecJMrcOD5lJvD+gXYeC
yZUuZPqHRevtPBrjtrfthicp666hE2SF8xVZ27sEfKUWQJXHrR3jOD9/dRYwkyCgObVYN60ccX/4
FHaYywA9vTtKVxCpLcwgvHpULjZ8mtwx0LZlUDs/MvCV+I9ft0t9eAsAJ3yVRkiY5EraqJS7dS4r
mMfduTolvbpOC8/yhnGxmtKWLTuwXqO1wzqlAXceG5LeQUgBtawn27/6tZp/hRg+caRoroWrv5Yv
vLQMzVseHKin/tMQvkisCJiXWrfnjTaJYsI4rAXtlj//vawqS0K5WeP1yRa4vv2WG7XU+YZQMZ9d
Pd/wcKrg5bsarO2Q0HRLFN313c+PNM+aigQPF7Rv1GfH/1e9PxS2Yysq/udxL6O4+YMY2LlalWju
tlAYNBa4Fp4o7TNXx0iDMzopAvqA7I3o9QTWDTfBj7mgV7du7Zdqd4LoyRvHiAK2KH4VNId4rPE2
01m0GOQBME79qZ/4uYcdj/TosnARZ6dj1q7sXQKll4qOXF4Xu4H763nM6M9dc11m4KVmfKF8G4U6
TlIFC91Yf1lhJxCkMTwN3T0oCetfUcpYagITiMmRNfimsEF2XBW86E4n7BZpxwGV0OnSi2aFjR1+
MTBRM1mAUd4MHT+O/PY8VN63wYCJVcv+iIhgkYTpo/n26fdZWM1ZGpOh53r1tASU1GKUquWX7n4l
v7rTPB6Q1q8zVPM301qhQUZVJlNaHnSO70It/c1/JmNMjxCVM7zpxcoIdQvaa5U88SPhX93BYtog
x/kmHwqbxkrqqOM6VzmSzOamBCRgOJRYNcYps2TpiU/5O1nJierQG1j02uYk/+paz4XNERssPHCm
X/kodvrieLKj/CY/IlBy+esm8S1inp1/MkaSppkze3PhxM0/hwJgAI24avlEbT8cKT6Snt/m0Lkk
fqzXtavW+yB3PwulE9PRJuz5KAaqu74bnGJP/5eZB/5xJpt+ga85kMgNvSXhaVM//EZHJv/leO58
irlBC1CYLgWrqgR59SHN8UO5qbpxITNkunMchpXY7U2iSg3DO08f4lCiUPAndcfVN6pccC8OF3ws
s8Rkw9Vx2NAfK7sMDXEljCmL19flfO0fa2CwuJMAiwkwJ9jOSZ8lCHqFf4e8lDyfklOgx6KFauwt
IOxkkVhh8r1Sd54eqy98i6tcKS2hBduoYkwKBJwJBsuHwU1RDAoLFJ7WHC08AlrwmSn+/rRQmO6g
nK/8Jcr2eT14Bhwm2sSFe+aDkEhbyDi3tM8Iq4DxFr/Lh14oxC/TjnOLDDcP1xDgasDla4LhaeZp
csTEDhipqTobGn+jIWtjV1M5+9+F3jJDi+nHO40/Q7K3NGSo5+XtXoeCP+JG5Q8ny1EAxQLlgpyi
TEJ36MioMF5b6m29Hh6CdkG+S1keGBQlMfQTtEbgm940SvXuF6YTWHkuEXrKUOQxwgefD+9CSPLM
hNROTnDzBfvhZFKQqtEg2AflQuWh4FJ1Cj1sojFG6vUEYwjm2fKis7eRwHA+kltshkoZz8Q8nH1r
AHOZCiH45ZhbyRORYGM26UmeWunFnlQ6yo3zD5gzhC7uRbDZED6CnN5Cv5OoWc80h+XejJ9c5ozX
mHmtkWULJOb+zee0mts2PV7SR5acR7lOICvnn7kODZ0jLIiaKY1OFD3nePv1dPkFCekOXuyX8t7h
MpuzpYbxa4H9B8eV1UFsg6D5/97imMIAuhsTirMaczPK/BtKCUMq9ebd07KMY0LueT8WtkMnRXTO
milWFaC9hzBVx1LT5ZW7tsdu+QCe/eSbuEIx7k8Emoui6zmRH5AEsxoobANaH/iGgGkbuO5pPCHa
rXxXmSYDEyjeQcZuiLvJF3bNpIjhLHuN+uqG+0PTmUetN7+MAV1M7pT8Ed0ApxoBnqqEDZUzil3L
up05tdpQyvT3yTZhinCVGBQMBbXlW9O/EuAkPHvg5uZTNeVarypcxgjRVL89WccBeR6+VOWgBEue
GYaR7BwmVuUZK3yjAbU+g6HnS2K7EnEAgMvh+9lQzZEQxaxCw8C2FnIX3gtTiqgEguMjzV6i36Bq
adMgGAMlCKVLj3+98claml/xPMhYJxTy6iJWbGfrdHbGgFIzK/v6hv9aaLggjvtgkWZDAqYxLTP+
b8JMe/2tD9ww2Ns2To7ckcboM9OAR5wSxUBhnKZJJ3BK4lqpIo6fRXuC9xN7p/yOiOaPFMLyZGNl
ssnjBvzcOztoRUl2TV0zp5a2k4y6nggt5whoTWLtQCiIInwfTo0/zbz/PTYSuqL3cvN97POdLXlz
MiRrnwNPz3aEu48SfsKd0Ce69tCUfZouHYkoPF8xJvNvVdpMzUi1pljDodyOlR7kCiqbaaBqNHAi
62bCCQlVEWyepqiSjQvfvgYiZJL5LgyR525KV5Jddz0V86oe1O44MLsKh9ac90N5Sdtic/0wuN9l
2NJF5D0Vv4h+ADjDd98aapShWqBYlhJk14bNK3RmzXVqqLLZ8dc1CXOSVysx+glmz+RDp/skz2ca
G+7+R39Cz2ikItr2/5DGeQevMI+LOREOdNTP2xT0UzKMF3fShb67xd0Joqs9iFkTyRlDS72HRxUl
tKjOCHf26JF+D1iQCUJV5CZUDCDNogl8zu1Ll4eYGI+W5UKyksVi75PF9Qrup4i2br2V62dMbK2u
dq0Qgz7qLijmdtRmMZW3I61Bea40458TnlsYWqx7AjFHDuD+aaI+wdJXCQb0rHymjrHyYBOJ6fZD
iIoD4JhOkfivQ1oQyt2XGpAzbZne9tPoPAp0yMxrV/Y0RN2+7ezpa2YrMToaX4PWQJgvuckhjeWH
lKOYdVMwcESD58W3MsynVzYSfKYVKgtvUdWQKRiPi0MJxAxY+yngDxfQYEAoaTEh9mP/mBmMHELw
qo0CTwb66vp31CGTCZ7RuYS4z4c8zHr+13DiXNB/bsLm5to81xblDUASrVmiFdfXhKTbE4Sb+r4n
8KJyC3gNGIsQ5sm63J/V0f8phcfrFLdT+RN/wutSf6zQTrzRiPohehETbLyCVciLeuR7X6KPwOJ+
MUfkhIrlzigVavin9HNYnt2G1Xj62DXhjbKaN2UFkGDT3ntA792U8OU3BZZIpaY2BdAk2thhIgHd
pMKHFnNUb8V3po5I0ok1woRMGQ+UMhRz+P0eMi8zfwq5Hg/edic0eLoA4271ls3wgwJfc+c/ASeW
KP/5VNdiUk23ZNUbWjOePrQfMvOdvGptElXPIWPLES9Ud1BTKTAPrHxmVA0m+7dboUsVv1T44Wq5
iM8jIg6BsP1E98rZcsfkB4BGyYuWkEVtYdNNdt/CDsgR56Zr8+N1juxA1wwWKOPip8OjOn07Jsht
E+82SQjw9Uh+2kb57QSq7O1ecj53VGSIhgVlGjPrAJuCrapOX4ZvYP/seeY7VWMWieOL1Rm3N31j
Ajuhb8OqwF3xtpo5wfMsy/MHgM5J7QZ8MJTyGfF/1KJ1Z+092QMQCz4F8BY38t4R9IQnx2I5Xt7Z
ISad6u7N21KFC/GMYFb3xS0u8FkL5w8IYf3+eC0pn5vaG1Kv/RurxpNv8B0BZvWxWYuY0+ZRvwEG
2VdQWVFbA39g6CrRgBeCMC0bhTYfGtUwRllKKl2UdBInx2NaPZ/BNZqRhaP6kHKtH3X4MMZNg8wc
AEMQHjb+H5/87PpWRT500xJ7awkpLgNf8KeMz5e+dOps8ZTgOOxU0wgzsN7WxUK047X+mw7vXABW
DW4yhhaZp/nGwfoH0w+2/SOmjPVkCijw6hFe4x2yEw1X4AsvMdAuccr5PkfWnjQlu4TLwjqVu5VP
FER/yg41T9LZnG5dH1+KhBklpvBazKtWgzoTsQQXxTLyR8+fIlggTAcfezejZreLywrOacCwSkg0
vF/UzjfEt5dJO0ISLY0T3lGeo5x+NcrqEEJ949IDtHOqQDOLc9oww/STa7MwmeuWxrcmUmPvXEZ9
VEagqe19J4TlrZDc1Bm5n5XP2uJAB2WPWBEUcwQt2jQLa5HuhdA3MRWdG62YF3WGo4b3gIFmEL5h
W+DmfkrUWde6EAzEWWh7kVm3lcVLCljDx/YQLTJ4kvmseSfVuOgdvoJk+CYrToOv8jeGMc6zvbkH
g5wlvOES5TD0op2rr0yMCm1kuWwaDQntTCg/ZVG9AeQfpm6WBO9n7tdm7YU9+Pa1034cpo9gIZSC
dKZCiukkYxXgcG8p4o+8YJzegzUB8C5+yFgwfgBgXZnYClAI24sXz53UjqpMThHrk+FO1Ypb1EWP
0rHjQZ4HU2v5P0XuUjtu7L1dsFb1F27nlLWgs9BeOgszdczKDbuTeNcoptEhPzYjEed7E1Q/vvQu
HDWTKsuBbNvwzTi9cci95Ljbdfjj88fA0H8SHFR6Y7nd5ttKwqhqZZKpcaLloCsXHHNF8EsMpk86
zvfkEAARR5q6PkW7qUwKsmIhtSfwZ6dP98sXxHeJD0F5qpfanwiEszS1RV6k34yRrN5iXQDAiNkA
7vLC6ZCx6DM1bU9un2rqVIXS+zcPxiwDTDPAUG0PydlcEBKqVaCE+ELoJGMIYwMqqImb0GX2CB1b
t/Y0Y0iX5xBNSYQXY3g7sQaTccj8dk82I7cyFJxz9tyoCTaNNkMG8G2ehoSDTuQ0D/tDtwS0HE59
oYHSUxAT5g8X1tZm9PiHKt/zq5XueiP3GCwGrjAbD+6aGCKwlLEr+8efLSeVOitr/LOb2b7nSeBY
R55by3ma4o23iryXorUnFHD2A1pZd3vN96/4lmjzDReRNBs/wNgbQrg5kUEeeQiEe3vnrLN7qka+
umhLKHgUGzGAvE0QLd2TUMFYnRx4etKxnk/CR9yPCSiBTnvtTaOSHyxMWm6sD96XieU4q5r4M+P4
KYlQDD/J5+Ctths4iptK+EoD73McZn1D1OwZUlBx8RoVvOv2bZSJqZXKpGVKWh0a3j6R6arJd/hA
Mwiq0ICVQZ2z5DXnfGHtdWoXVC6l575Dr32UkWCsSU03B8dnEbzSapZZyxGe2P47KWZnnkrc/kw6
OdgDvy4MF8ByiIBP5Hz5ccQSTsM9SSFOP/PVz8ndO775lGyHq3T3YJ2PSgETlmYws62ploWKxoQ7
wuHllWi/iEZIOlM9W3fZ+SVwU2iNh5MLWhfJIXzydDlGfF7MbQ77d+dyqdZVLIGzX/SpjCRVMa0T
T6IIV9wxr8Aabmb81Ovz5PWY0R2oXPnz+pajhm92gJEPBiKMlsP4I7mcJdOpFM6bhSNzExmtdvok
27bpupHoWyySH23/H5VqsiHKiOQoVrYcT9byPNHOHV9ePvFOz85GflugHDMO1Q2wEtn5WCkh4D5m
cUwzGwlx5CExH44rYnMRIyvTLHFmoEBaCNltSsGifO9lhT8pTqtq33GVUhEfN+GtbPphS5z2kNa2
qNuXH1OZ2Ttd8FO4TNbvoJYKoYI73slb1H3haaTVw76j8yMZrZMDFjc+3CfaW14IM8iiEX2/dGsB
RRFnbI2602qbCayamWlmK8DTAV9yehlihhoEWI8QIAf3vHJ6NflGfHzKvzACbchdk2ByG08bhY1n
cWtAfm1k76HGM3RSvYTjJD/UJGezNCfa2pjZjLx9smwhlssjVWeEKniuUdYTGBN3EShlQDey8hc9
8bVlzPm/1vl1sh5ToxDbEUXaC1y4OoLyBBEfZaacMiWQE0CN502c79Ksm2mrHeqbw5TJqgEPfAXB
xxJ37Sxw1eILEr7vmZO6AHhW7/LupJncycmCh5ibcoM6Ertwr9MOUPDHDrXMNy6ZkDKdcA8OGoOy
6eKNhQJyBCpph25ipeqpg0/SFZEh11Yr8Msi9AMPtkY8YCtVjLjIueFLkTtLEHvMml8Wl9HCUAb8
OU0rMsqvBQPwtbABolEIAbFJxCQuHWfs/ijL0EK0GUly7cXuKA6cNlMTgBnMYLW6rfQdR5z5+3CM
7MS1maXKulAGeZCceC0EJgDz7oOfJt5bFGtHiE9me/+8Z+zpn4ydsRcuU1E02gwfrIHPw2Dle/p/
0bgTfhR2hjM1Dnuy67TRXHn84t/Eqh6AXIQtkJy8zprCpufodTGC2D9pSgKOfB38R6KTDkRWGG4t
GqFAKqwlAszERqW7b5d/Ny8Jgv3lh3rB25ty5gAIlHnps+qURVg/a5CeuWzDWrN2eVVFRRQiGeZS
aAY4Kz1gsyX3oRWmN5XsasaSZaO/ToOFLZMA9fNdFEpOr/XtR1hOtTQLNealzMCd4uRVNK6HJy/6
HzMB6FlhJeKP3GxKtydkD7gFlTg23c6c+mFu4eP8Mbdw6b60Lw2a2f0u060heqETC0rl1ndQD8iw
3fkc00S1rfqRx9PKZjY3JGAhxFMESCf8dnuZP1ZBcoYyyh73zPmYlcF/r1jMIrExUQmABXAWgFFd
QOlkan2bfL8vHudG2zK80LzNZbGvnMJ9eB891Acs9QEqcwV+l1cDc5UUMPMvZ2iEAB1BH538SaXc
arroLpIAS6jOaWVimK37uU/eL+lcV3TuRdALkZ157HEPhWlZST2Q5NX9ftcULiZGHqRN7m/IhB7s
ebFg17BJXQBEjlprNV9TuznS4a9ifvaTetCPm1u+KOKRosZPhtKmV63fdD9baCQfz4TDIrcHpQnD
PEuvGiuQlFvN2cFOblWNa/oKQ2YKo88RZyRkyFzi8gN9mm2YAhGIHAsUk2z4TrhuQCLegyU+z8/8
kJIq8cv4wNJIBo6ry2E4W53z6vnsC+wMJD7+dGH38Gkoi4yrsAgK1cS9oxb6+pdmBlZBwFu+HTFQ
+w2zt6OIBIjGk1CIqDtX3B+CeUNZOpo801zHr/c0Hvy6GNq7W6ENBLxF4pvkitkg+7TZbMl2l2nn
9IbZP4gO5zAsGbF5zQ/OTvxGVxMzWQ09W13gUUfe/S4m/EShW5n7/15xOJft8st74xy63uJDJrGq
axZP0+yQTWjojVbc/B3tTgmeTMkArbt3t/XfMYhiV8h6586YN7O3rYhQh5Y3KkzAozQHdJTJA/9+
5g93yVYJO+whhMPSKbzVonRQJt1hH9H4H0G3cle/XaLazVJLB7/FWQW96fMrDcbcU7D9su5hoW9Y
GLeMu3/HGxFjCcD7Lu3J+dOJP99DIsnjJ3zyaXknnzksKzQDGdTzRdDAPP8foH4hqShH8aPJCFT9
FDe77XEuFFzw0u4euqDHqLW4f6+zl9fzj3t/cMdMHF3KvnPtCLFibiHjVN3Y/O/JSyj43+eqWVHM
q1IvbRZ7xPL99C9e+EZ/H7dcxaK2mKwT7O/3aOm4pajpxDrpQrfLKZsM6LCRq8tYArqasUKs/Des
ZqMDlbkqhFNCwVoLXkjko+7QMNl3xA5MpLYwZywc+zELuZwgv7SDnKUVzrnuAoSl1T+CnFoRFRTz
8VHM32t+NUh9zWwCEAkzHT/o4T49CmsCn1nWK6Jx2ZLI20Lbfk22Lhj3jSmfP5jDu5zMXIFyRu8c
SFLWPCaWq4ljPM4rrGcbQb+Nc0d9080Dix85AURLsmfy9qqTe6Bd0kKAPayfJj6uIbVVeNog9rwx
oZIIAnYZHgMSMoeNAqkSMeutoOImkX7ZOfiTPCFoFnD0la6y8ftq8ytsjETg2AvD0X1x/ZWptG0j
n+Ujs0ylJY1NHZCGjr00gtM4QZtlmgQHAeun/iAMpgsPeLTUn+3MnVYd+BHPujk2nhY5R09/hwSp
Ccp/yvbzaB3IIz/7AJmlrzXanhIERzvECuFpde9tEz0NOOf9ncK9hIm9FtfSwvVaUghEKugb6jgx
nvcw1yICVM7nMa7KCuSurAeEcxidCbU5/Bf7Y2h5xQRH4dBB0xfJcYeX6j+tetncqAbWzgfm8qv4
5+B3NYhhLo1h7dEu3F58T3+CzmCWmUWznFfe07D528ndXn0OEMtNKRs9Z7lH5VgkM3EEPtMbMpob
xJ2tUNOXfp9ND1A9kxsI4sQoWNUNg8eOhHXwu3gGawBtkiYdwPKwK10KuPsoX1lMNX3SDgsPO6JK
03klY2Vqzuy4QxySewElkxntIe3RP0960TGHXCOBhjmgRJjJZXJu5FJyJLWEaOStKw/4a7/e8lOF
wx2F2HNUICq1Hs+VORoro0zipnvFdd8vDFKj5ZVnd3y/Fj81i9AxLvl/wHJPIxPyEMWw2EK72fSh
B8c/R4/CbPD8st6uWi4x6XYTCljHtrMQTmne5Vi+LZVQh84qtFriO24xWScyE70SU5bfKOQcoZsq
mxyeh+928GUujAuPuLJaZNDG53ZeCqOaFuSdNUQFlhjEp4BZOTxfaDIaX462CA6J7g2qEMhy5hmr
nKFPAkOMTmm/EHVHTTjbHQ+3gLpqz2KnDvbVJbmP6B63AGrhn6akDcj92LlkA+IC/UOiqmXkHSMU
GjfbZM4XlFg4y96lCSxgSKg9FndaE/R5qyMPc0dhINdh+WSs1SLBRDTdRHEK9ZBFTAUatt6H6SAC
p4ieI9KH9knXVLYrDWqs0nfzHSjsrvlGuZTsWKRDcorwdT5AcdNtevP0VipYs0WZYS41PhGZbLe9
tjrieasPT65hKwklXloXqqGMl73qVa5UCm28QTihE/mawU2YyQUiZpn5jlCPRTqD9OMm8W4h5nre
1pem07C12s3zMgxkD9qBGNobUPadhFyj5VuFTpbMELtQsZSbrnZt14NqOxKZSs09Tgz0t9uZUQ39
t3yT4q4Em4PN/g1w/zKwsjCod5ypU4VDJYQyee3HvL++llcDsMyLxW9RWALfl7eFFPe+ca0gLAoz
rAVMpy3GXh/13IZM0b0SF1t/HfpKhDYwAHTDhIram0zsOSzV5oEuyPtEsp2xV7RmKqFYmA9/Ep3g
ewwg50VewNPM2GkUFGcAaDbXL8o9xZXPPE9LHOldfkxYVpBiFpaU8eumiULjpcOuuyV9rXD4wGyh
XQhG1BrFy9YS2GeOCYyRpZYtc93V+oj02iFGnlRB0TxBTdN3/4aDKDGwURSsygdLDhQxdjCxtioC
QqssvDSmt6qCknlmxYdzh6mQO+geupwbmfLiNW46b9pcgQiEKI6JQVCe/Du7Rzc5fpLSwDFTPxhx
YajRlRd3Ul/pSWwhu/FdUnosLc+5M5bGMiYJyQQ83jzpM8pQCfyrx4gTk6PmN6JvdEr3ZPIo4YtX
5Ka3Z2Z7puAAY+Fq4/KVxE2HYxB7gAMG8cs62V4SMgJ7h/QKjShrFf8w2UdJahjB1pBVfRt1PKiv
sZHhVeaQiE6JzBp/WJt60MQBF6pgV/ylLLkP4K/Obiy/HdB8IjD8e3PmvgjrPuYzIZII7M8P5YmH
Q0oebG3Q32dRPapnh/8ZlQgD0GaIKe4gvPQbhKi5Ej42A9EM42m36UtqIzaPOPBHqKIoa5FGnsgS
ZIDhZiK2tDeFfRw1kB2ufFP5LEtG343K9StGgZ8I4U9aGHKxhjaGCanlw8zOtIUke5vofZM//Qs4
bYG9K8ionQSWdITIPH0Tp1AvKlzOvfMJ/H6DVbZ5rGZqYwFvxcf6G3nLQzuX4wkx3HTCjs97KSqi
dX62GQSEzIQRxrIj59vvQZN/Qy0Ubp5W7fieI0art9VbGPb61BqKFAb3h5L1EFWd/BHR21GINVaM
TkMTmxx1ka1nyqvXPHB0BE7dxYNxmBhpe7O7wmN6pMZtob5DSTmrkMYmf3/Vt02qpmeBo8FJvmcJ
kD3xPmXFZTQfBlG2h5PWzKeCF1HFFIlkuHc74M3EDv+8TPnyPd7tJt42zNnrdgBuRR+EeCvQQJIh
wyCNG1/9Qo3kCxkYuzineS7/Exfm0Kl03VR8iQ8ABjOChyWlTNn6B9LwUE83J2FkDgzwfvYzb4r0
zH0dHhxQDj9rfKjs3gGEK/8yWWaZ5LT0GzEExSec95MjIdu16zBeJBSX4cZs6AJ4VjGJF9dI5BBi
XN6Q7UxHV4U0xaK5AeO4ZYoAKr4piFKX2A5V83ONvkDq5aSOeKHDpy0A2jHmN+EuUxCSDwkItEqf
mTL8Vvm69YP/684UXlAtyVM+u69APwz3QvHe+djhiKJ+vUIzXq4ufeA0pQJ6STNcIESYmvrd1pP7
XlpIRnYZ7wr66rKqTKblDAjq4hV5wBe7r2GB0hKFv2Pw5igQ7hIRg7g13aszR1xLC3zl7c2IJE2X
BYGFO4JE9bCAY8PhFBQo4rdoTvDFk5CAoxbhjW6wN4ofz93H6MCaeI+swBl96BIS3pVI1dEExn1E
MCWDB1Ud3YTURyQ2phAIZx+RGr23XoUoqalJOrtAYTK3bqErMkQn0ogfnkaybcoy+orCqj5ThqH+
UUPW5xoy7Z0Wc/RR+h7H4gisNHkZQ7m+u1aaPbeoyPdjhZGClUgbJbuOrYgagMeBrd4snEVRuwZS
lVVy1iJVezJUes/dDjBH+zcwh2wQvGREXB/obra58mOWLR5EvbWJIkni54cIKHehfnfGS5NpIFtT
nb3RsrmtJEtFatRQMun4ACkNSIhsGTpaMHk20RI8aRSr/XmfcMKFFZ8I+PE0JqoPpezOojI0LCHT
fCNzHwtIoxQrE9QrqVxqrB8muw4SiLldJtYwvdNb0R9+ORiVvXoPu8Yeoa/quBMOkLCmJh3ICL8B
f9L1uBq5hFFAyJ//Yi26D1A0GwntQZEaDO5898SplzpqaplS8F4UcyQSPSI929bjTNZx75SEVAD+
AUvWt27/hl8Zg20iDUiBDnE2vUOy2K4ZSd6mvxk6G2vZzDgjcVqwbpdA9tnD5oZqkX0vawIAGkh0
K/eAJ3DEOX/U7Y0wxD442h5Q36F/FBVGLxhAR7kkdSVKJJx8DmWtsiIXeAp7KZ67dL9L4//Lzdtp
JALrt7Crzs86Pat7OrEbNcWPuH2KmteWdGmGRKFn4ZEp6INUcTlLtmmMkq9Cp/Q3FHhkNwtFqhf9
rb2L+1O85Fv3/xc4WRVBOAsTtBHuq8+7+WSdlZg6BHuVO6ptMZ3Oe64tjIhURCD+/1x4CuShRBHk
gE+SU59V7YfiwYoQ2GFpSrAI1v9zE5Rv8WjQlCWKacbcVqfoWsbzOylohq05KQ5b3BR7Z4g5VnKW
4ZOuVOJ8kKmJbKHrvefJ5CjHDFAlB/yLO+yl/fY2KlN+E7szUJR9mMx6cEhziy6l4kBE0eBLh979
Yn7vj+C2BmhLB/yMPKJOb8IOG8VPmFn5zRueImf8EL97/847za8ZILC4v3aUgIQO9CzBsFEddWhP
ynn+V8uU99BVjFTXboG1iz27w+WSpgdCAanqayEpK18X+TPZ5JQwP8Lb9WPwra+Goh5yBR5iN9dp
zxu4CY1yH0lkrOfEzy1kKwZ+noRFLgsb28c7jVU7WbeHgs28Zzx4dJBacAEMhgpWKonkpG+RrTD2
jcfLfYCkqUWw5RY/Uhy+V5DL17c92E+QRCD5yGiyT+7ZJtukXR7voS26vGYj+69V2nHrSFdJmyGU
/9hntn/gm4NR2YQhJpKRcRvrgMnzsDZSIpJCcweeROuMr/isXSI1+2XkMLqfYRRAH6R1jJ+DKbY4
bP24NJAyJius8dsyj2jGNtLP1UpT2jTbi9Q9rXDzbn+dgUKjP1ZDBN5+hp8dHfHPULRfkVyoApbE
QyP5ylwOTE2cJBY/gVgT1WnEiYHmci2/ojLxkGMlJ4p1tgwi9DQCVNzUCDrRdirT01r3io/GX35q
uudrOKFhi2DrKXeHE24Mv1/DRto5QKN8cocfZfKPOcxMfS2MUBUZSGsVkylt1Fa3zJuao91sKIIU
BO4lO5q08+8A2O2MKW9MXZBkofSoK5ZXSX9zKCWIj9j+n7E4aE4PhEegcViOyicTD0rsmHfnRGL/
EvqMCEMyGX4xgVDYa7mJ2qifKyYbNRgW46mplOR/Qhg2PQRnYE3gqsmIkU0YtzQgSBT1RHE39XKZ
jt4cp27nQOxFxZ9rsgzvrhY99pZ08Ozau9mxUYOdGdZVLYRXqC9JOPQmqbounIC4jXA/1qT0KMU2
aYdyeCSCv/zmskMZnAFATd+yusUf6Vnq8+ElxqeYajF27fjpYbEa4Yo27X7iFVo/ep01/KfXvMw4
mHqaZPokCGr0TBxWvupsQRryGpuhgc8yI9tKo78DeXgCBzZ4pY+fE/0y3A8EQvfH1oLqmgkaVswJ
DwdNp0meq3Kk9shIhLXEuPs6vJtwh9TV9CZfyaeCI4A//MHa/9QCsaxNlA+UugKlAchzQeso2qzM
0BGBnMPZKoZYNC+tRMdUBDHbvWlyvptqsqlONeQXtthtWD6HbzE8MSrzaexgRQc9MLIQjE3ZT8MY
dv0uJbmJKDRRyQiKVEbg+3MlyXHEWGt0DqpJKQBjjzXNc76OGDG2AXu1HaSnActP147yQ01RL9N+
T1vwbSlUFoBYU3VJ1Rzlj0qQa4lurBjCreoWvnb1/eTH/siOKAl65BCgsaUrtkFnR3wmqawBSpUx
tDMkTqoyWSKuwNZihzH5s89jUxCUdTybzzhop5rK3VHIyw3jnllgBrkIgCUv8XlxDKPwIS/3Es8s
iLMxv2t6SbSjZ2BUGNo9BiZud0p2rD5xJGQYFQzlVmPrAnBeOxUh6n1kEaS+ib8OSdu1u2iUnHc2
aUtQVyIh5sieTt8N/zr15qft7gwy7hWF5bLV9UePJw+SYzx2a1J5q/nZte9mjMBQd6FlLOWTtnvJ
29L6ktrLnD+EklEck3PSBMUWpHrPyiGElr+UKMUXGFXRavnxL7d0G2hxZxNHxhngxjNdfuBXNpxh
EjcZae7j3jMzs+ugZ8GU1GRCWXgfSC6UWYQ+wSuh/CzIX0jX/5zToqKKdU7n99stuPjTZLbLv7Xe
OGc2p1B8iS4sHX1HAfyrxetrcZqeS1l8ZZ3ZzuCQYsegx0Q4N9QYUUr2mToDwm2CaBa6uNGenUFJ
SQKibsUrk8+C4wyi+BlX90QnkV7Rb5l80ddBw1axTEdnGUesGWlSBTCR/SffV5N6oqAS2vp+RRji
LtsATYsKRweGZclqgK1k5Ncooh4NXDwDnDs+yZrv2mgKAC2pP/GhrLU/CJE/I8IHchLOGclLAx+q
/8UqDqXa8ZYY1x+OpkwjHhylB97kRRuAnbBrr+tHmsFoe/cwZ/YJ5tQmEkR+vL1jppAqg8mNtfAo
opOBS93mEt4wqfbCArM8NIcvWMN2xqTMk3Y33hmhzvlkc2XdMt/G3Ion2v5IuBt5crHOFQ8DDRNg
8JbyXS6UjI26JdGQiV9PNoOraYdTj1bq0T+flDwv8SnzlbldPwpbTUfrFjOjMCaXX5rubaQylNuH
+qFw9j7LjLsW3BjsnXy1iXBr8GcQv4hMMvKSvyzlOY0R06o2EfGPUDtlgl0N8hkLqmcfqy+dfUKP
WYuOotawOoNGAXx6cF8vVRtVNMJ7l4nwgTJjkfmGsDGletcUYeevqdNF0uXofZkEPLo87GyH9PR3
DtganVsWCyO/eYXVMPQBqWJ9xzZp0QLVUmkcdbUdRR5io2EH0hCRNlARm8B9Vl0J6+ref5MV/t/G
9PMtHwC70XhVR08yuDEbaoFWhlllJE5KLAkX6tlxBM5FP6WNmocP2wDNJmKFpw632mmG6Q40Jm2F
cT+PeDAlKP8BNPGFjPkmotn7hemKSSpE+v3GpW2fhxcP97uGvra8PwMCiK722zd7vRa4XmBda37r
7jIG95YUHbYVOyJ30dKel9iibQkkAt6Xe/Hg19s6bZaOBoKCPhmXtjMJYh+hZ/C9w3QwUADUXm0R
tDmQ4gYfDJgRq8pF8cGqMIIeIQvdyy9PN6Qk6u2HAYD+LAq42FcNkuqiiUbyNU/kgLMZfhR/8Nmw
CgvgnqS7oouK6Fx/m4sbGtlAsI7M3Wbcb7kaUzoRBNhy4TOgE8MsL5GvIBvP6mQlOsSZXkEI5UP6
9u+AP+LoyHHBGTub6cS6k8bqH+bDOMzy8+czlR8nkXhj9vN9JNhfcbZDzOkmwApSUVVAshZtBAhT
cno1m6k26eMKWZJ3vGHB3EsECGnRgO7kBzIalnVuNfKLzb2w/OU6uk9oNPAvbu1FN0EYsTgEe358
RGeuWleK6jSQE9EmdyZO0geaVFuBl5aVo4c+ch0MY3iwoZPYgAXCBSATYti9qdXtJiywMhl9aAG9
McMJFF46ve3Y9miYj/ZHqQNn5xxHtLl2ak7bwcdHruo/dHd6PQO/GQqHy4dX3EPGE4WgNNDnetmC
sOjnmql30+ngwi/vleNueaAoqA/YYsM+Hec+xsODcPXBm7V4bwdeRgIKVlsdvncMtvlOg8rzYGQH
jci7hLyp/fo2ifA9rQIyUE7qpPx+BxQ6v30VLtg8BLxNfK/yDVSL1HGQQnJgg+pj5Lk1OeUVVnIs
Q+vCUAZAPi8QxTM+9KBS4OLw3FF8u8KsCo5UmU/k7VA/5728jFONf1XoNrf8IeoTSCCXa5sq3mxw
x9madqoVg+wxKAnAyqxoa1aQCuS3nbJflirMYzQsczSBAGQ2wwU2fX87CsN3kxlwQky4zAhSe0TS
CiVa/BiPyenEO/MkKwzhOhq5jrpCs5wRz7UiJMqA9Uo9iU/rdcwwTe8CCTNTxYS2IlJu/82PBy6+
Vi0gLFuR2fOUWlMsG+s7OoqECwqjyFrvK9hQFK0JDAt8nu5htaO5MpP05V+a3DXQ22Nnfpkdr3sm
oJ7v2l9V3B1u6F8Xik/2vyR+pj9XX8W48cBBS61KWXE5mfSPW6180jD++optIxWPTIfG1PjL1jhy
GIDksCt03/nZWXksEXLZ3UJBHBIr00NRcHcL0z6SciANll2A3v5t0sGdHwYMxeWoEIBFeEtfS9n2
MHkK2TojS8y4uHjvdut///j9LMscephcoBWT8q6bnx7WUyUmLMXTkp0K4pNpEg9amEFmYhxkejUf
mzFo+Kc8yv0KuMxCfjZcpoaF8Qs0RnQyYTDyGDrBptiav8idVaA30n4S2fxxLnYjOHrhLhWrk9iA
MbENHmjL/aHgbZHiKIOUhJ2eLAOBjEL42P2zRKkZTo1aHg9dPW13lKQjzHKjZVOactKfRn5VU2mk
AC8MnHx0Xndsd1o31ax2qU9g5FmEI8hvSWMiYPEezjMogWjOiCD692ap6Fh370HNvx44YFE0+VW7
EbojAwdUHncKidOXW91ArFLKG7DmYOifo8ZllI8RnSlDSXYLWtYdufZCyIMKclk+tovU87/35KOS
330iHoGUDkD6Rov1F8PIqrEZvK7mCMyCfFv4BRqN+QDvWHgO9HXi/+dWHBAensjvC3SBoEZmJwI/
uIPLk22cZcw68SYbViaJC4GLskGCWOwyMnxFH7WSwG0LhCqJy2WCJrQcByH9wdl4TGuYc1zn+5GN
hj3SXJMcdUXl4ZBn3E14CGhqcd91bu1yWQiG3fXbzRjpEeuXkl81IYBRscXwnazLaaPUwyUuaG1m
+RJPONQI4E+O3jYjA5Hmb4LOiYfOdbxpBHXyTMSx87L0bJXjR7pLqKTkIPvqxS2lfiMsKKmz7E3y
+KJiASHsKpRHNJOwT33dMOm/IjUxwUyOqc73R8cVOGtaoTnFQw98/TODz8jWA1bglH+az+B+KrtZ
EQ2sOr3D+NVXucdsUMaUgggz9/XV70DG1sWUM/HQcIz8gqi7iVEc5tJ++/e6KiSj9oZTca4HFMMe
BbvnE1XnZhfadJH3hVMPliPjp/oeuN43Vj1zxtVQ6DaV2+3bXPstO0rUyEwOTfhqXM3gJhM4cmoZ
51RmLlBp5kzT47VfPoCHJy0BdBqxbtY4gTNM1ZCopZ8U0vX/mlmHrTA44yUEvu0meq/eL8jdEoIG
OTDXcs35NqdhQ3c3thK/0NIvt5ZGS8qanNuKwlGJS8K38RJU2+p0ULmGX061aOJ7kX+MkNKT1ZrI
cAUQvXKgNcA0pu0m18P2ndTHYvltor5jLZE7X5BAEm5Pjo9BDsqfDqSUaNuwOBTUFjOWcDjC7GQc
JYXkcS4CbiEwe9cN4MXtYLYNFGLIkDiNvyLh34IIusWan3zawKwtKcDju6CzYLCm2p7nOBawgc77
ZTzwNkarRERVk6IGEhSvJlr+uQstD1qXtkbB/CJWH6XmTnWKPXeAdW2CTR0pjbm+WDWGgZTZDSCN
UlCnYtEXF8cq5/Xk99M2G9xMZi+hs0y8uACCTX7A2SwwZproxtqgLXHgMI6uGcz5kC5Rd4xur9O2
7AQe0j/G514bk5aG4A3ULoikhCLjKleLYYLOAahcwDVVjS/s6mJH2aFXyDvl+Pzdr2q9ChFLh6rC
R/+FOuR6dyBcsMPJ+NUalBNtpAfXlBjrfCooc5iLD/HjATCrAAEZQYGHDZawLEm8Xvs7ciUKeTRV
Oc4uZ92/KB+h/fCIgFE8V//Mmv7RjxY5xPqER41THhu4iByx3VdoL2ohXQtpMov8ky4DCJ61rNp0
Io1XaIxM7hISGkccGJZKO/K/O3ooRicxZay/Wcrv2P06Ue/zOfMstxqWLQOr0XIBdOtlml62dvMK
GCezlUjdkQ6oOC+wUdqIEGqhc3seT9CY0YZ2aKExOjK0q3iYAVwQBDDhRIKsB1ne/5D2XjO0YzF9
wAKp3T0IevWGNjpdHDZRBHQNIfK2jrRwUo1opqAuUnoNARVy8f0u7cVcYWC9WO/nNrkS10aDcIdB
/1oBKy91VQJwJtWWmAVWBdJMPDreS5BWkgJ2wcdeyQ7R44hqmUBtHTV8ZIViiMJlYB7FaO4lKpCX
eI8HYQ7NJS5kpSmXLIwFt+k21UGCR+7Yup6HWfjb0mD82NJNR/AOYsmmOScQsZal1RgA7cexN9/F
gXEfOHL98nKjbSkitj9BDxbGUTauDUJC0adT+DfgvCKWvdwavT9c4vlspdxPuGwc+WkxlcETe9fK
+dx4FOBvuq4VJqjq/8ol2M8SY/QutFrqSmZOAcb0HVtX1ekJ522bomPfCh0HnzesaXh3eddbKOpC
0ggF/XsmB9R6XwQA2rfcAOyBSX90gUiL+UGMtYJNfExk0v0ZKiFqnQQNG58Gs2xE9xl86LC07Kiy
XGqngjhkMlA6lSIS2W8sbXUdsmrKKYAqacx4cKyeSEbyI595NxHU56o6Ro5MpbKttB4dtTztymnh
JhYBJklQimMfg+46Ffg6h+nfybEHJqBhZmXafQgahgMnZZLSWM40FdM70yY3uRH2+vGbWoq3K/Pu
KX7WNjpVxnySn+RZwbHvzcuIwfdI7ewUvQBMax58HM7k/Rscd8Oe9d7GgR6Ehm826dwc1Yq2ke9u
zkgL5uHw9BP+TY35KcIBBjiJsuRHDS2ed23AxPiBR1v0G8cAnEoPPuCGrmqO+cb/Ki+3Q61Ivqib
8CXdYwidvmOb8Ecpfc/lidjJh1KWrqytaK+kxeAJ/D8V15/7NnkRViryAyk9UDbCtvNkqPJur+kl
tZJDdEUI13VXs5NGIPoGyAmRF/7fMfYBHa/IrOQQlDW1S7quSr3XxG31s0UO1d5wj+4EpjM9AUt6
SliJoBRBtjhefy0yNBpJBOCLQg8Phc6sEHgHNSdEP8ZL9K6iE2NmVBkII1ouUrDbKFXijF+UaX81
WmmC48scE7eSO3AvNIygxyUxzLlxXYyXshbuWOA62nak+5VApOkt3FUkSqiNsLA6ZaiZrEO4XE5e
MN6K9uuL0lOwVpEcd+/NL+lLph38RfiYJ+pQ9ASiKrHAJ3Wk102xpedHPWk361amFamykU8sxBJO
ZhYA1IEYYuCjayraf5JZeGTChelqZzDe1y+36YAvDG4u1oly/QdXhz5ieWzPIqNq36/vaQnA0unF
F2t/C5+SPSA3bZBMAm0q5GCx0VG04HK5Pb3FnjwY1lAT1LpHudxNcRwKjBPTsVjCFwCQb7RO1rmO
K9PvgJXD/5nu88Q8+Xmn0okDColSBIrLj8OFp+7nqjlQsKRRYfhGrbP0U4VNgBiFTyHJMvwOHUEi
6p2gCiq9u5hyH7s0wH8DiEFx1z1TxxEKm9Cow5Igsqmbsl+0wHEVZP3/FAQt1rUmE3KNKe1oHTSl
1cJxd74JNK1fDimMzMqzdNnj7+qBPy14xb+kN6Klhd+6dFepxjyqCXgnR8CX0B8O+hlSx99PnBb5
Gqo0tc8JXfTFQM/wsu/6Ggp/53nYN//okUAzrPU17wK9gPWtyNQX0TMfejzL9HsXPvZtRndnD5zE
eM791CpvovIY+j+TyKmJp/wpRs8y/2gkopWmTM2LxQKQSKWVHCtXqo+YvikBj2MVG/O61YzypCJ5
H31kI4gdWLFY6X2lzOKO2KMPOc2PHHJp7dmILdyu0naR4JogXq8b/HEKO+zIMlWNLTC02RIRCcPI
Pzs3IQyiRNaMqXZT1CVe2vsxDDbbTlm2YRZx0ji3NCufuAWBIVPcWS8U18gvnKYJySi/hKnXfxDo
/+cStu8MycBjk6idHzLlHbGGEFYUGms+3Bi9NwFU5E91VMDaVdx+gW2kfp39Wtq2S15Q2T9MonnZ
R8kToWDMvDsgEF+JmhfGM1hXBkxJg81Zh2qYAuAY1uzNolNwRf7IQ+32g1BWuoubMoVH0z5kCwSH
foJUkpfBcgyXDZWOnsPLTFoEot6va+XWikxhJsUh0zxuM8s2cyt/NvYgt26+XkF2K84fR5E69ANH
CyYSFlot71NsH+oPmpHWgw3X/KiK3/CI10JTM+tH/OBz0jnU82qUQ6KlfJKod5D6hEtJBn34lH61
zb2in9HG2brHu2m6R4RutSO5w5oRwBQ+wHPJcOrUNsA6Tb9SsydcrvaEj3eD+shaNK/dXJ1g0doZ
a+1j73yHWOgVVIDR1rwc4azs4Q2e8O0Sm0QUjFy5vmhuJHt+1KQLHnp2OpHsgmEHA/72ZdDOIzcZ
05gy8knKYGojjV456UY1lIvjqRhRjOXs7fWCKT0RLUOCE/w/4RBW0eTXrKSf0NefaSjB+0sbQ8x2
bOanYbAUpVSDscL18oV8UYti/FWk8GONolyO5+YuSVeeYXcGh8V2eXJyP7Tq9nTFN++BriG6TLzv
nL2yQ3jczY+7Wsv3dmJgG9uGwjVunhHlxjc+uPJ2AEPLbt/7beYbiwNCUcjbGjBx7NzqrQFpgpKl
Zu/MUV94A1d0vK34KYw0BxzJxba3yakBjTi++8gUWgE1NDtXhELrXU7iy3/W77CbsaWIzcexu1QX
2vXJKFhqX/6fDOV/Foeurp18M6nQArxnivoH6XP+byjw1byYFwpisqZ2w4bNYpBFDV5ClXMoj9Jv
ozDWpRPxb3gskGa+FSJOgFumIsAuFVC6I7coxUkg5PTfmyXVCkgtTY/Fg4r4t44Q8G3/ShrSH606
xHTc0wgVYklQZSZnI6MCgfpVZZY0F7a1STFbfO81b+nqpajKDvtNUJAUaNqUTiTLL4LCrZUZbBrX
NAb1WGPtJhirEZ9hVlhFLtrBWQIB5Yc0v+vTBxasj/iG0wl9HlfZSPW2RXQoPqVyfMShub6U6EDD
SfVnxF9+6q/KPn4R8GJajhhyOj9T9qABmbV/XgrYateO9tRTcWty26G/YNKB/b2Lzmv/5ubEbS6K
FiTBLRvrdkv7w1x+fjYW0G+PBJnCi540YpD9zC5Q2jYiseVaRsZO7fdl8LIkIFaSn90/ndnP34ba
dWeuIRynKp6/cF2xHeWewKT9YrDlLfvpbgJ1VOiNrtTcFS2RUU/4+dceb19BQ8BLutRr7Q7i+YBU
Ch2LBpUJJxwoRM9IGwB+0llXDXjAjwjK5nWN98pAZxGclPwC56Q79cSAeO/mjQexHVsPLxe9y1dk
96KyIchDZ/5XsyKJInUmhAEaXYKD1wjqV5xOnxz7pnJal0qugZXqiShTKd4zvE4oTFrbanNKkWMs
pNzr5mfok9oADqlcdU5IExaJ5PmiMErpdhz9lsweS3ZQeeAcBHNhO2CJfrMCLD4CLHLP7mXW3F9S
Bwx3hvplI5Z/8WBfHDm9HytERS4Jwgq1uP0/xqAFHsjBufqk8rbeYRioZJcG5eYG63KHGXK7tTkK
MHOpP/hmNfNfyjQvwY7jxdEdI2zg8tdL7Wjxwj433encq05GGcgq9kDUO/nNoqmMVVH1P+c0i93M
y0Ze1kNIgyeT2fNADk9F6WZL7oS7y5sq+A6mL1PwkGW+82MpIi24bsnsEd8aEeop+/CZsL+n5ePz
fIFE2d+Z57ft5eGu0mf0YvaFmU6dko3oCmU2dlnAgt4sMLdJeOT7Pr3h4OO/h+131cKgRShP6HbU
Ib3T8UrF+/Fzh1+yIHUoUMzpnw/HRzQYwt7NPWRM7MOsFXxOWsdGFd3SYOSOoUhJ8Ldiykn+jH+X
/IoAmiwFMbMgnsdoec4Sr6enRiQW2P2WD9B2DiBdaQPP2giagwNJLytMKgqJnD1Y1AR0nLmkYM+L
Qwq3+gFZHJWCqPoPCb4vlwJo4U6AUPENgQMlurAS2qkgkcc0OQLiTVW2sp2YTU6UePv70PzYIOIX
+xB9c/gXtUKqsaL30ZMCGNiWfa4IgBkb1H1a4cSM0oYPc0F7feG6RuYfZowvGAH+M6JMFexAUn9i
vC9fqjmu12GEK5lywnWMhqeYtfH8Pd/0R7xJld74wJUUUrWn2u/L1vYEEhTmEmK0XqZrbp6Ql851
HvX5Tyi5DVU8T3CxjDcRBDlM3gKOFzp1ArlP+f3jg4yD4SAaxPQABAgjeHysKBg772IyTi9tuiYv
Q9HAbELMtORJMpudbq9n+8C9ScbghU/ISvAMAYRocUkbGjzDODrujotGXr4BHjZJJWWMOWGY+o4w
JG9YOHm2YA65SBryO3XztcUWuuRiFDfdv/9pYHMGKsRKiqabwZApQqzKABZ7yNAlHjB6pDe+tai2
WtPGAVdyYjusg04RpEwgibxZfTwMez9ybe58YpIgN5UjENlqB2HNap1mFpV0nDFtRu3uvb484nrH
9NRSJyJArqPTWBnHrEOpwWef5enxfqfdhpNdy2/geA1UAa1ZPtWWY7CIe9tXlgOI80oe8FFrvuaL
eAEhez6LcRRtfagR6o8e5UuY0ljkF+Klf58pvO4RZ3Yf1dv/2+LFtqhZG+joDHcwbZBYAkuLEt/V
FM+7PTn8eEGT16N88mHyt24zDjD+Qb2yqsu1N+Fp0Up6cSPSbMs8eZmufvpa0l1U7oQ4zY0aVph3
CdEH/fNQZP8slfccy5ka5avvR349cZSqrByB/UO0rXJAlS3IT3eBWJCqYJlCzNfPq1EVkgh93VoK
cWrf6KI+QSdj5klMk3ZU5Tf5TU81YzCM2Efzc6qVnCyTHsAUrrj8vqVkZobU6LIaP4TXD5q/3dH8
fW6rjN2T2tILWVeSl4buXN8Lx44qpIXBXFAX7ZbLRHOaDFtZ4fuo+ci4xV7STDQJhf33qaVF/0Dy
Xe2IAXzyq9kZ3ttBLiuBNglBe6/fO0WIQq7E/PXxNZ6+q7imboZqyIhig8TzsocW0eisSe/fwFGy
Fh8ImFWZZwMec6tusteo7gBS8R/xI+fC2vWXNZVCU/gfNMcS0PIoHTltjIa8FSutDpDkXqThxlLN
9LyD4GSvUCN1xksYz/Qo3bCf5zZs6TCsSH73yd7zzsK+n2vnIftIVc/E38tSQZdNNBtWbh/sBFJT
ZZ0NbmkiqiJHf7doJ/+5cdGsN+5Ugnfe1KPRWOVM8kcE6ibRyqmU4Wmk4/TGg+wup9+a4Phv11cY
pT4TPmX+UzUqsIA3v7q0uU/Qc6GN/qsbRYd4EYg4rupS9WRQRm3geG1d9/nJ1Z6QQJupsHPd2k4M
+kBPVLsCnEaQ4HedZHgTybx9YyfAAfPamF/87lEtbNflpnHuYzttQlIOnI2uDBnL3Nz/YED2Wdhk
OnJi8KV707foL39R0atBfnVEaK0AgmxNXOlDA8cklfGSw7fQrRPAN77DkA6y+GmpsBKLIhIV17ky
HEJYUGPXAvnW5aPuVgI2LPDNi7WLHyg+YJvvD4ZLZm3OuDrjTxmvwGq1d7dsIOKB+Hhqy/2h1QRK
Nvku0TmtPm2WgIE2BRIXI36HlW8MMESGQydUm8HahtZP/uA/VPhhYLXzjS+LOmS9McCTEOxPMQc+
IZbAJ1f1TdWs3bT9zdiREpJjyroZ8hbBoL4Hq0i/Rl/9au1ZjCKcktqBCmIPc9U3UPxeG9kouNIg
niKggxzyQgy1Wz6CodO7K7exh5DcbY+11PUv9pJk2ufGR6P+tvc/2TYJwiXX8GiLJ/lXhmIyKHsF
hQXbnP1h9MdbFPKbUAXNtEVAzOL8G4+8m4EcNUDBvF7aQp17qIjd6htFp8pZ0ZnhPWqkfEjUBRB2
cLIYyMuL3tmrH3eQrQTDmS/uj4OLVMnXKhdtcIh4Nc4OlLEYt8J1o2RBi7+l7U8KAcvM2ZVLbgRx
Pk2e+w6gx1OZdGELZA65byaTV24IjGbAH7VNVzs6/Gmb9jUreq4QfzdZrO5Ux+iC4Uv5N/Vbe8Dy
c+d+IwA6LE8rWOYLTvB/AmmIC8+7HE0VfxioFCx8w684WcAz+nTtey9NGTsTJmc00Me4sm9rEf4e
mkbym5tzN8U3qe5wN739lbMUbgHwVC1Mn36UI0PwD51KnbjlADtbWiVUko2Hg1Rbq5rGe4ZEH27C
o+gwat+hyZmYZpOd3aqWUv1fqViPDyEgsvXeYQ7p5eNqR67RwvEt5mVQaXI7omw/y2qSXfUuOljN
uwhct24+CBImJo3wmQzDgWthdh0/tyxE5sqCSKiYcASdx98F6BbsuTL8EzySgJHdsEmDBLetxnga
PG4q6mPW8ipuSYIWu+JzcXs+S8KsONgJCwUdPtv10FpDnsDOzLOPcOP6N9/5sb7nyH5/r3BPhgXy
KhqdVsajdUu+7wFnLb9xEd3Mpr5EX9pXzp/5wIoy6XQy/mXFlaZPPkpyttEKBVXlQwGUgcQRxQ4H
d33HEiL1P4spICLxwvYikT+sXLoTSnYdSMtfqeZmFPU4dabYXzXwA0DEDOarFxVBAyO/ACuq1tOo
TuyG+3zTbCyFX5K0sv+gvSGAZoM7lUNZioX0IGf0V/9UVmaYE8l86rO/6TStVSrR2KymI2koTppw
yOq3j/mCsn3MuRAYb/LUTHQGJ8BkoebYqS4uYBS9KL9zU8mtY7brE/CeLtY50yfj8jamFOmqev+m
uhs0uk6s1X8DNp4bXLBJDlRf06pNMvZ4QYL0EXbiQGHrh2Ruwk/k3n4LS5pBojMu9/hXhjmL2JdX
qJJMhqVf8LKkNABeYbQMOTxLghU9aPMGcTCAWaaoSfdWHA0q39ot03BFvABcgc+JyKJDk+nZ2H8X
7UOBvhlJjDumOQIy08eRPhZ7vjlGaNlts1zrHyPAYUqGWU2UmaP1WFcMqlSO2SCd6dhclrRUNLle
ibdORz1q7VDauGyDLOe4sQCyL6MKBX5TXPQMibop6lY2iWt8hi50f8CgS+fwcy59rKkpJyuFQGu2
N54VRRo/i4CE80qBWNq+KIEJxkz1bVhDVhNvh7qCSikbn9+OJ5Se50z6uGaXZU2tI6R++o6X36GJ
Rk4aol7COP1UqrgcolzyeTOR1dIACXh/FlaplNZlVa1yuiUN6F+PCSlTrAZnaz0LikzU/LBqx9K4
y+nwbpXRJqOaQueAqPiPi24Y+qBvGldwgVgzq4puEpjmC8XnEbLZ0PzVgYN/kXoMQNrXu1rMxOrR
eWcAGz4ElnsQ7hSJOsdL7PSW1YpDx+r/BpuJ8EucE4h+8hoeQjSrjKEFnvrIyPp0f0xD0XJayPFH
sVeFhtHTQSwCQBgkVTw8bBPvQiLbazehO7Ey7FZpN/AcH9GWcZ1r6Y1kXalktThmPoSeT8ATtBse
66lff9F+uhLaSjvaomE5eBJXIUitfvZDzKZ6/WPdR0hXoylgQet9TJ9Im0+fne3rxP4sa8/gDCjt
jLKWzjjBaQthxZubhBuDN6EQgxNUuSjypvsIo+A3XTAwYYGdFvvqBna2Hz4DIJoIZSH6ylQr//rW
X6HtGi/q5vFq5uJVMuMzZsmy9TQu0tZhNsQtBKfnLRq4d2C2W74rPPQQoLqO9skfWN7lkHxpETBW
Q+8uohUzWVR2s93Y05MQftkYHlmY+h3KzVFUKka3w4h/Q55QJdvq+xq8Vs8N+6TSZxhneEw2JwcY
NpsttzD5zKudhIoSrhiYglV++FmbU82LbrREnz/rfXW5Y2M5Ct68hGYS3Cg5SO8C2Lfzn2muq65A
ChWU4c95HlpSVskbe3+p++543HuxZ1fgCKeFCB2F/DLhLoNB7cp5+kOHGcI4P2wMfL87IMSpayg1
IKK7XdVP1q2pFN10W5hNFQpZ+2rAwvloLi2wSq3e+9+G6UkkqmbsI7LziZkFA2N9CAb2fuhtyAJc
1dCYJ5eNQj4NpfmHe7S6hk0lwbZ7OWCRCYnyG8Wegud7dhbpTzuYROY8x/NGbvYTU7+4tON6ZOJz
8/oJZMo90XSpW4qb6KYkvajhDnaELpTSFYsvO2411nr0c1uWkYEjF0PPdsk6nD4V2ygLKNVlONO4
p6vzOtSt0snOJXABi9CFa12M3OK8GmSgJWze56ibClcE/AF7KHTzp2DL73yAR6v9jVXn1PF2+0uZ
BP9a1LAgxes7BE3e4IrhCu+t3Rq0U7STbdpVnxEqc3Jru9m2RDidXyK8A+gWd6bfFGfBPXQDuKhY
EOatGbyyEHXH2kfOVCCDneH94p/Gyq11r+r9WlwIZR0+28dR6J1LDUFw60aiU+m2xfj4U0BQ1h00
pYnsGsDN3s6mWMnuNTfUXS0DOdstXxzcUjxZG2nKrW5feXQcvDUTNzahjJQnQoe29HVHUL2mEnDn
02TRqVWdUCwWd7Wuta8khNRyvoQ0w2noR8+MnnQz2L88rwPQWS/uKXpc5JPYUAJhtCpVTfVn43+A
zJLEzHbCjX8711FtGpkyu8FRclnyg/o5CxlLrKeYZvbm35nQgEbJNNd2NQFkOySj7c9RcyIF/xR8
nrMQ5ObFTLafV0qeOogxK6Q+4iHbB9+CcW4SNQsJmvpQPLPSEaAoQ5n5d/JiHgaENHov9XR7qeHW
2OCNBaKIEWnu4ohlnGReY8i/tWFcB94K2IZzRW1EpRw/YDiGMjDLOU02uAVkvBCxwtVNoedsIPeV
4yR+ZAstQrwu+dSz+C8DzplTsgz8SeaJjtYtpuqvgzVXG709YZ5MYinM7QFgPNjRBF7yKr6qKWcr
+6WfvEyKwnX/9PoQFfNUgSKcjRR+pfC3UqnRaC7+SdZ7n/szp5nE/tOyfGwtlsb9qNpqNzSIl/jr
0t5igd4ST6XxMOI+dxGnaoZsDGm2XJtiBdQtjPgR/SDXATcVpGJrlk7t4ZyfD3Z/Y1mXrI74qQlR
k0zQI3wMOMTqnyN9mLSZk2k9SE4oE7bpOs7GPPmu1OcRetbSv3hs5rMnW2bpqIdSHn2va4PIiVL8
pMqaFKJcGlpzk5YmUvyEdafA3XUpmI+xGvazamflx8zpZZHdNuvWJ4gUhHC5+vaZchnGnYBomHGw
zPKUljA/JLAHb2d7FwOud+AaDbgRMlm5wO2h7Zp+OgJoW3j4mqD2cHQ09cD3BWmqFiNQenEVi9D1
tYZn1n177LMqqlwoauG1FWq8FlOG7/ixBzW0HyyxRaPgQrPpMcs1yEBXuJ2ySEK/hQNSOXwmJKx5
YR+B5V7G03Hi5ig+1NGg6URrs5n8maXEazPnZzNi2xgiJhRKfPJ+ulSXfTBS4bxX474VTmxy81k+
6iiRlYke4hPzYevt5wvOk8fRtOOgz8OGbG0GNs/2nJWMfSKgNChw+YcxMyDJa/cCrfjEZQV+XEdR
0lEyr4Ba8ll4aJos807AO8F/I389wIKs6ooxdHxU7nntoNKSWdtFgysbypScUWPahrJqIg+qIxy4
EyTwHan57wwTLig7pSPygehqlTU4lNqM5kWqO6pQTvbhumGFZFadyU4SlhNpBgL9dkkrvc7mpKC6
5c9OeHNazNjl7VciBGMJivqYLaawrPs9DKZdxaUkWQxBo28VNMLVFV66HOjuRo3OavlQTrmAqmL/
q3NoA8AszCFTeOlwojVCoNmC1hWe7DWQFGQSAX3z9AFJDm7TtXhV2aUthMEqkcSUdSuHeCbeRCJR
KX+1GYWLvUhS2dg7UuGMbeYYETg1skZbuFyaOU94qHWgTusGES2PU8G3/UvB5tZ7bymssoL9iGz4
xWZu4njrZRrLPx6OTf6zgiG67VIJDjbYEsElw39+5fMMNZGEm6XB7TWnUTgYA2HXE4YFIHxSj0yE
BuVHuOIkWsSSrI1pDQIe69dF44NuRb1HfPWxStdZyDr/cTfZEpGeIAtYRJP7So8Y+VE6t3HNFUZE
Epw3yq6Atjir/RH/xc7nltDAyCuCV4z2mTDpatU06j8WSCjvgJ3jwtCESpGuBceZPYdrihVnAgOf
wpFueOOr0qtYPFliSjyBJOtvbDIqi7ETANzxnlWlNP2IYlQNT5OvEv2dY9CP/VXH4O0hyRvhmUIR
M8f7WX/6rVBMyqNUQcMq2fZgwgZuWwW62u0G7dKoalWE6AkZp35dBuIGw5pttLOFR/mWCJcpG+4m
pdA2z1jy/nlBx8MRSgCCReMx6SwMcA8GDrdYoffVXsLo6SgoU7PP9NuoWGuMHwB/GN9Atek8Rxnv
NnUtN8YAFU0NKhqfxsJVAU0fTmGnwPVQk653wvhp/SIBwJOAXr+wPPo7Watdux+mCrCNzwRbMnfC
UJ9qkMHxzpqJLtWzUSZ7KDxdcpyqHKpYpqUl6ICWPEQ7nruiMYyKb0JjkYeuK2f1VhOQx5mla3af
iCRV+rbhI1FPtSmN3/D253akMC7CXj8WeYWAHA58VPkuA64nrH9qZgOKuPF+sBNuwkH9b6lt8KxN
y6F5PgAT7jjFnrBF16VHZI9q0feY7QHgLPp3r0i/q/jlK4xmqx9iVUMFNNHl+KvABFrf082OXEfN
6p2h0j6Cbm0xbPsLRDa/sreGWuzh2Xd7JxAm5g6rU7h7MoY7dCK55+QoFD8C1aY9Xp9jaGR7cxjI
EcuXxERcELI5FG6KaoD2cyuuoznSRA0KVsb6uS7OW+pgc0IVRrZIxFN6diwUWTx2KIvsLaVUffvD
UdD47t8oJHbkeI8xaENE+8g6e+xf8qhXjamj+cq0tkq+JD2K3NBcgIwsROZPaAqyi5pbdr4fvmX4
9id+9nLKqB8lpoy0JxRJfVu/AXXY1JDvb+Ez5HlodkCZ3H07bUawrUy0/4yIqlBtT5bxV0DoJbOR
KIwtzhqCHIRENQsBNtUbd5e3iCVEI3Ys3LelmXEGczkjN7x/7VkqjPpEwnfkOlXSSOgS5fn57K5J
RMDeHbWT9/lGMSKZ80Xgeki41VO98nq8BIfxR30yQtE5NRdNIDB9vddlkZydKu/O2bYRKQCGWDZB
FskfRfjiGqcBx6wcA9Au1iF4EzUwU1RcE/wEXqF3QKfLWEiGQ+lP3CyCXWXDXIxwSzDsph5+ZdlU
yMOmaJp76HOF4IiAPFx9YbDAGkzs/o577z/uHi9n5CPA99HmQEdX5QfaaoyOSu6RizpjC4oPLY9x
q/nkM0pPPbU2N6mgnOBtWcj5l9noAI77WFYrCCnyALmJyodRzhKdl+CfuCk8phIEarlWl/wkGJ3C
PFEb2CA0SCMc5O6pI0atuwL3uDiup6XfDTueiEJEk7Q4OtQmmCjsn3lxMirCwY937fdblR4v3WDW
wMap/8ZfP9+C48tDf4Lw5q3fhYjicZFXeXUXPjLmo9qVGWxDg1xMeu278C4dm4x6t4f9JXHQ15XQ
8DRq4SMnoPnyVd/1gsyIh/3Jv51HFFnXPm6qdisSUFyO64hPWTam0HdPEbpFHbUJuhzg8E4G78zO
xruj6501eEZzzQroRARlWHoSA8bXj7adXQIwXM1ZBstk43vPra/0+Dol1D65jqElKcqe6yT7ZvgO
kMH8/vRDWmEug32soRi9HReLm4x3o9D7vKVOGv6eE0jMqGdyxo5c/YINzeKkvNYV+aMZ6vICpNHJ
aygSyGvJdnDPQjERcjjUgVhufvM1kX7ORyUPRmG2rIWwBlQpGPjHQ+HXVfbnZfX7F8VyHFZgzS+E
kq+N/qDxIi5L/Ioaa7b6oomqmAgq9TRft6/LImetvTJoFslE5Ufy8giRe/iMK+gFKKafgOZ51rwo
sEjbtMXf2RjAdr/LVBKZB72/PQ4Kv1bvB1dBXO0KQeOzDIIf1SBp7BCViXCpzAZvp0zQWHqwWUf1
VDImVdnpZI5/OiVYDawJDQIaJyDjEBALhoRHA2E0l/Vv1dohHtcZh1zxwME07tY7+KAYq03+Lydk
i3z+y6gVU2iQy26AZ3EwW4RmyZveucHVbrMt6nxdmXl6IO5Q0OZNkJhuCEpnETB5MTITCDzh47+l
zRqhQnb1JmDcseAlY3oc8DY1ICrgNVJkPUM0EmNSDXk/ZZ8BBH2TP7fhDMTmO73SrI3T7HwdtMYo
8wpEUMWA8zwzLkEPuS1mcR9QFHOtrv+FAzy+fmmKTYNqUbNUzYa9B6v3YXSZHsm8TjFbilUYb+ge
l3hRO9Um6NXZn4PWAjm5BeIsML2Pgow6A9qFUTCth8PTcNh+BokoOE3NomhijyfLk+n+YT/2SKvC
OZpWWJtxsnhgB3R5xqavWpCf//RxKj0AXfv4loSPcXIJEZ2uhjSRVPlESrDFKI1ZsKhqfQccxJKL
km7B2T5MNUveBPk+VMogGiwVIFh3D1pHGpUuefiAVnaUeWurrsYMuJRIsTn20yAg//hZ1oLAG4oq
q7FtTJT2WaAMeM8UTyLMP42j8v/5x/0Moba++aG4QQL5nGy0+uZ8iRlpoDqkQPg4KgQJraILAc65
Y/dUFpzWMWM8vc6rZbXc03UiGvgkGqAc33bZsSM8rfPn7H/JSfTvzVBMM6GgnFJ7IUf0aIiXJJRe
S4VCIAuEc25DtIdNbdxR35y/kuxgAvRmc2d+1cPApBTI0Y41IlgmmTlEBcISo3JK/HcmH0wMGZMs
a7yY/Qq3PCXGeCzr9jpdphEcSEbQY+1Au00x03kMvgPyFOyypScw4zCL6E8vmm6sTFgsepM/JkTw
0knPbky9y5MtsKaLiRPF1SLOP/3ZrXDrwFm9l9ya5K1evkhzPr+xBNgjHi0ypYNMylHzPeIgwOq5
7pf2cdwJeTU3xNtbr3b6TBl1iSi0RRCAz6zlaL7O4pyIsWrIerMnz/omse76ectXdchQneXOZDi/
/T/p87azgE+yKEiuKizLo1V0vwJWPG7Gc3g+eWMR6/VqekbLv7rmsdwX6ytp+ROv8uT1xM37fMyu
WYD6OlwAwadux7+OpYaoRbLQ4HPcCX/CC9xZIVXrBku5QivwvaycS4v+7pP28us45Tq5MSuz5t2N
HJ4sZmUsbfasGE7CBCcu/5+N11VRqkNxP2YQOfUTfIJnH1DGpIPjmyuKGQxLKuaesjVTDYzEZSKL
89EjwxLjCPByB0C5+7lrONCaBWj+yu2wsjPpvaVLWjany1b3sHteeMbBJmEf0D8C1JhyOjLaKC3Q
9uwzKo7SyikMrKb9ajT40LY/8XvgEGvANfcxAskt8BGZHcuupdL8feS/QPnQV46pCqlyittnMfhs
T1B7QhzTkzR6yOZSAa7WWaCeD20p+ZNFqjPHK5WGUY7im35kp0O+UglEs7Kd7o/Ir5mhml2py7ia
NB89DcWQW3kPZ5mCon1RdZ/XZO/qJRCQ6FC+PrH90DTCr9ngEUK9RwFcScbgPi2tltyodnRxEzok
rFbJ02VkQkazfe+VxmIMTrV9egsfpdrDIUU1hYSjECEhTBdBFeW4SGZzTFNbg0mcSFatNW7ZJ3K4
yT5psQApkvBXllZjf72YruleoQ0l55BuWJHssAvcDqH+opRRW8kf/FV5uUVeqpQKedlmbB7oHvSK
k12m9sBX1QGriGS7cyKRqndVZg/rwUTwhKqjb6ADNlV7dznBLi0UDMMgTs+PGn05NYPH1/mthOrB
9AamVuTr6A29lGZCxSz1kFCgHMlK9+Eu+UKxxJVEEEEHPovdjWBVO4btu8GMFN+Tia+/oPskq94Z
L8VywH37VTylyPA8hd9aHa8OOT0RW89JNC55uedy6qPdZ1EDS60Ufb1XEG4pne0TrhuuWBH5zcHb
9XcmVIS5lhZpWPapo0nfC+4K2WORsk5qpZXqy85wHWsgKSYyByj2PYypLK+QpiaGEAHXvaXNN4my
ElNCipAs+NuMJL6cCXPKWdRTXL21/soznX8WINqUSVE//S+NsMwzRghfSnQjgT0TFu9Iqc0pe96+
BoOA53A8W1WyvOQVyIs1GnCefaEIllDec4w9reyRwM6sy0YVDxJPt6x5gWntxQwvcpCpr5WipYFg
2fdk7mZymbX28EUZAnFm8pJf9fTkXcGMCiB5NsAR9nCVReG5otGIdFLWJq4Dl9ga30YAfej2aw7u
C0DNXZq+7lyvot6BDTdWxnb4/3nJ27M15QsSnGN5j0jJSbXJjQi/wYPYecSGQNnb0kJOIcg6WYtR
zHBi0CXyNhIatuK9FVx7a+/LhgeGRUiu3Qi+4ZjDj4Uk3UnchBCAg4pO/fYBeZMLG3WGUWaTfEAb
prgM2nuOEdOhW2mCNYaLOrt/DiGvQx6QUmjGgKVQvvYKqFECD2zg3Ksp1Xu092Eel/K077ePYNSQ
o+1/HJxF7BoY95thalBy4GqW/B8DnQNbOCzdJR6zlEaVvJIgs5qJ3q0EOGEqpzoLjeDDoVUf2C9I
ZrplBLdNYsCLM1V44zCBniRQnFFA2ugMh6dOeuAAk4UgeO9Sl3ff2GfAIO6e2zlUaEUeFZQxwKp7
OCV1BZd75vHg9tm5mfPLTs6CFN/gdUXgZoHzjLYuVjdTy7GeAR5fd/x+dF/IyC9mYi4h7sn5of34
c8Bx9B5ti+SbwPHB/vmuUFMRFvOKzXJzdtTk8uTmVBX/fVcVjL2rKFANGA3RHJ4PtQyvd9wsrS7W
N+8AFRvfezvpEvpqYG6zQ43KmqsivvgT8Idya3j9N88Qxf8UV2hbXPAq+Tr5Cw82Mtlu1dnEAJ5D
uTXlYP/i80XZ+cjCShVWLkSCoqPfM7NkxvGqOavcv+7/58hhW7aBbXzt1y5ZA+NF2UvOXuRyyhj8
YCdTXhCPGyZ+eLZPiVstfwgDHerlG5LaNHViYV4dln165azt8OIq7M4lrfkLCuUPpOFO3FWHv0k+
zFOqAfPmu8OI3dEY8JKIfpW/iEsInVLEE82sesrxscZOJvUPmPPHMQgsms1FNVuvqzeUn3SJst+d
haNkHpx+qPHfQM91Q+x7tSH4HbhDV9gb5LnVf5inoPx0qtne02AoXptJ5tjrFauuPMZvcJEVt0tn
wHtO9wdYUU6EaAlelYBxKpQ/GcAgw8bDK6uSGrHPtvVZGrIv1JfKPU6z2bbDllHnn96XgQD54+fE
S10ZupHpX1s7h+alWNcJR4+AUgeD/pAfNKDfFcnimDy9AtK8PMvt6pPTUjKJoV0WGrNDl8XWc7Ef
10tVLtC+uzrOIaY4xIi4ECi3gIIKDJoWGYFmi+31LQfW85GYem/V5zF/AGDXAlmrV6eY56ZYed0S
HXOaZxZnJ2YXV3PQ4X9FBuwZ391coUsQ7A/pvIDrYZ6krGWgZC0+BhH7mApKIDI8weWXkAUN8af6
ED7cJsLS3px3chq+v5/J0EtQiq2BCIGOE/gaovgBS23dETIx2Iepk6w+ZmFRFzOnFDQItYF2K+Ma
aEgww+VTMd0hJXRPEbsxWZ+eolYEQXJOeplOLreJpXQgcTLTWX7vACpYfRr2H/X2+1+yciXBNhkz
8ht9K1b8PAP5sM1ZKvWIwCJAydZgQJOUTMlfhWMvvXhNHm2v00A9iCpH6F2CR7ThBX0FlVjuTPuf
4Seme06ozelXCe8fiyXIuv35t6bh3dGx9v952f+mbrH+PFLePTZL7uPMMaGWhlRbFEOykZmMIUQf
gDjxluPKjwFRshqtoph7GfZISRKJ/ibMb70ajaqjBtdA3K4ShUHeqKSwHyie9drCG154LjfXBPJN
Ye01VxwgoowDUY7yBB2ZWxGXbsy3e1isci4ySoQPmASFHlWZ0FBMFYCjt/gKji6QSkGJWPs5YCef
13h0IZsNwoK2OWkJ+45yvxSugygN5rTSBL3xUeZvh75t8Xj2jI+F+oIb95Pwi/WKvQcaYH71nkPC
GcYzB9mJkPMmDbBGoTHsiCHCH5bDc2Vp5b/9rYTPNDoJypVNrSojcce1Jxt2Ok5ahUpnlr3UfncP
oVPA0V9UFjCT+hhWTQgC7/MTMIn/EGM1naMBuZr52zeSNk9ux1rQF0fkCZCrfVALCnUIYskb3xUO
BRbMlIP14ZhpYRnlM/2amPbd3ddw8uidwX+J2U43JNePSPTv7PnMAddWYlu0BDxSXBueKnIB9lA7
Y123lA5j5dUC9t6HoYzmM831C7FkMFcx/ETW8MsOE5TlaTTkWo9/yLKl40Y0FaDLemvMLWAQMvvJ
9vTHJn6+LCIvt2YNtT1r6PFerjXVdCf/99KNnffwQaH9kCnuvBSlxcHmIJwDgmv2IHNrOLdQH2yN
NWonj3fIxq3/NwdCoRKlUl8/Ky4Y8m9DT1QyrWcDMnACQqqdaiGeR+SJ90UNdTGbeL6CKIorqLp4
TLYIKOOznGcARn9dF/X23PaT5UFDmn6p1jMFSnVxfzvfB4BEX05bh/KF6c5ydsLvWW1MRJJy929H
Zz929SCTQ54B+62ZlJ73Huh8Vc4nl/CNJ+NG2pErXDMhdbsNjRyq2zYm4iNyk17GBHuOYfCEqHzQ
gmILdXjPMsSNx53MZIl3EPnscNz/7QgXZX671ppOF/3CaYFypJDBxPJ5KC8js0K6+mYqcrJQir7i
mcKP1vTpYAz+5BfONl12hzL4wRq9JZR8Ld2SMVaG7lA57dcPYkmCjejN/An4jJ//LCuSxwTqzLsV
d+OA8+06j7cb2MhA1PYlZE6ub+eLdzaZrJQ3HdbQNTmiTgNy0AYLB4lUe8TotN6ijdxjOG6XUaXs
lxgHj/bWiO0QZKuEh2svr1PHofNLt/3pWRNW9H3GQtM2MyMudsQLEOaa8mL/GyaPVcz9qRrmNOoI
gzSt/BMadWZloe/DE8oh8rIkVlV4LAHuYgq5G3tWVZYo7h0ivYpftMpSVU3kxS/YccpwjJBv1SdA
1Z2VC9FJgLPmimy9XsfobwpVpfuaMSLpsX1uorDk/qh0q1r2yV9WfPWCk76xcqp1Ph6jsaORJYWh
wpOPLX6OHhGBEOimVDjP77p45tuChFkEp0NfxMTng0ESm95omhJR2feme/Vy3uztW0XDRvWfMExP
McdldmiydDK390mQHQXxBYWQf9xgaeD3f/wis07QXt2dALhnUpmPRR8AKTGKO3i1xSpIL2x7Zd/Z
p4C+FOvyk+ZfLYBSIwlRXEoL8AUUga+PCZhtzzcC+hT3CZipnbN42PIrw++iYKty/GvFaJtV+UUK
T00p+wXpmqysrL+JOB2pkdG5YQ/cQJirq7WqLb/IshcvMkG9mef4FZox2Kx+0lR5sqNKNZCCdYGn
miUN329JCDKblfx3SgkvGUrl+E5R7tm9HqfOWEe3JdGncjVZ1EcQHdkszDyXVIzDNdLgAg1+fqia
tj0bBbMoZ7EyAc8zMAqH0xaepFlBApnM3ittD/Zg0byh7X4aqv6CG9+UJNp1ZVij2/Fv1RCZmgCT
W78BA5k4UsSsyyJegA3KL3WtL9fdZP932ik4c6omHU52zAdsm2fsPsS6zywm270gqEucqRxPTKn9
Jlo+Lm5encJAssw1ISfMWUnAoPtu+pc5delg0oFMJr1pxtgloOPPA9SnyNa7EsEll0e3yFfaXzdQ
6A9t6vOfHxBjkfFelxmHwpe65aadtjxbtz/BwxjS1Xyh+nQrULOm+WG/fkJow388CgxqWVX56AWV
FKVxNo8VgC12/ff6Qmy8njz9kTfCenspzaQR1JUKhXUrWbhdvRYDs3Lx8Y7TwS/LjQZnDVDGvDCx
fVupsVi9FSXVAnKNN7VFCYjjXDtZyfqR1nL1++RWDDljKWAJo/QZgd5IWFRoNV9TonsKEmcimZTA
Kzsp7JmOfftgNXuXHeLe1DjLgIPgPYy+2AW577MKjCKe8ogfUv8KehPrnRsCYdR8UX8vEXCs3nqv
q/vzOcyYiHSpfd71ADfE+WJWVVtcpzl1ZO15pyq6syyQKAQ51K09nqnLNn6ei2fk5z1Y1iAEp+81
P94I6c9Gd3kxyGHd9j5b2RN+aWBnKvuWLF77rwhSr7naZZglMITgRrubqP2sIJKKWtmhzq8zWSAy
7hll7jHY1MvcFj7WvjcqNoThyAfeQ8GsIobi5cdxRg3K6SbJSDqg3+qXDOHy2b5UtvgbYKcZUhVe
lwWkZqkPZmlebo2tPxSmSOuBqOhx8XWhYETszO3zo4QhpgHnvqcS4up+EXmtlfAP/cKj+Q37eLPl
4CaWoUWtwFT/mcq8pOK01u/BEpbC+LYxOK1imK8aFN4GzAb4kPjXPAVfCqpz/MKnZ1whXl5XuxL7
jrn3VZ2+AKzUedu/NA/EqLME7aHkE+L4HwEfJVqli6w2UXNacon9ZFQVmZ6ahIGJ2nhBrl1U8JXv
SnE5pZsjKwwCdhArIbX8wNt0WhF+R3BJdQrIEB6MNlPEPZztnigXaAGKou9SQ9oeov/e0W6H2EsH
d3Y82rcuaUtnMQH7johN1qzr4jM50MfV9Xyrvu8oAZ+4AIPzrL8q7eI/j4ykf3fGRivuzR57pLCs
glPToLohnAGGjXnMrg8w20Rb5tDd8wlwIpeBlAmMCLBNvKDdNsIZcYsG/C+0jivx4Vm9WqsCrSSY
g9TcssbAjK81sUaggPd9Kbd2OJfLmIEwablVsqbkHpVEk1dgLAx5YH6jXQMNaZkucSFA8n9c+DOc
j7jCfs5agOskd9GnWJLEcCeJ5QrlwhSKRzlZI4NmyEte3tvvr6YZEe0uOcki6V7Im23px9g75JD5
fz2euoKlpD7YD0anyNHExwTirFn1xu7mvW/jhEA80ptR0Xtttv4lDrTyvPGeCbx7T34GQkox9kLt
yXG2xiKyV5DrL5gL02gOSsf3paAdhamBu48ELeVOimgmZmEUFGbM7y0SP1udXlr4yiLCmnKlueLC
zu9xUppqQBa3O0d/wOm92tAgtJq4smWf0PL7UslmrJ5Jc8NRpl+EUIdpd/d3jF/AJL7YLR4m8P6U
iQg4TXTSNORgIriePg/cAd+XpxoDiF+0WCj7yIIALFfxW9xc9itp+V/kHcjMXElhma7XIr8qmzJY
zzV9u2oBt3maGmgZ3XwLR3FTf9lab26cEfHDeD7UySLtWfpZKpwnoRoNPukwKVj65nOAskuw07WR
YMP4+muP/ljxEbhZPGvoQST3xGiWmwDfcv9sJVee2DvULhWSgRABZ4amoXrSD97cbZRt+AL/YXKv
HrmQfK5gcU8tSbZ66WgCOTGcSa0XigLuVVJTnXPhoMSLUR5OH/lg6PteplXqxdcgnLU9VxttSQgC
6pmMgQ4yQEBeJ3+WnHJZD18mYYmDJdQyZ4lB9DV4Y1zoAlyygc3Ne/xIWWMGBdSli0yQQ00fFP/Z
K+uNXoa/60cJMujYTLiZoczhP2050iIbrme0opj0u1YvPHLqmWCGMibDABXoD/rZ/v4hi+ZuEuJA
Ba3k/U2X8YkoAcfF20LehODPICx8mjz5yFfPXzsNv/GhVPTWguQIw9sgDEZYY49/HPijjWFVz0s6
QhxPy9p54+pXSafkx11kANbkZLkTj/zf1vkM1HQmrimnBD4cjSnZGE6Ekj3tySNO3IcCcF/bkuDe
QBf6aNSXrPcEzlQ00PClUPlukth1XX0cXFBW5Jg0EhTXN+bJT+Uzq1wC7Gg6pkURxVJjy86/mQfe
oMg/KZvztnvp3qsbgUS7hfh15tTkPUONk/8Xj8uv9lA2a1tCc+RC6xSArnO47LQ52izS0mgqawyd
XQftoux317kgj+UqZv6NObHeRUo7r9A7jqb+nRfrtEAVyD85ugIhU/O1POJW+l0j7MRdKo1gG7pD
9e6/fCMFeFfxJYE/rDEf0u1rF1NTe5/gi5JWPNtD5FDyBRIgBggecLqn1rGvmCscYRNpgGvaAWNp
ppShg+PnY7TRMlCMzkJukScaHm/kJF4wkNd0F6mThbTh0GvNXI2dAZ1RnEM7uzv3nJ1my7dkmXqv
EtwyBvRgPCsUlVfaXdREJdgJLZE7fl0rZr395Lj6m7Cqji0jAKtixWouQpjuIJrODUtCrDhKpEfG
RVQEFfMhq1HGFNXI1Q1I4jcrtM5TBb6KB77nEasYTbcXdpazaN31hLBmFMzENtIPmVXXG761wPfb
yAE8XtNYiigUnRp6vjsJC1DfApV8iWlscnua41mbE/30GrYAvFN9zMQc2JmUk68z2C18eNQ5n/rz
xN1XkN39mgHj+r2Q/YKYxCCFpe1uvPi1+05tCkepkzoa1X4U6CrCznD+N243QtVbVhcybHzGKHHQ
5dRSTbVEqI1yRhk18w27eGKod6vS9op6p/8yyVcWIugdlEZUiHdlqHbVNgoNqCXMke5Araa+HjK+
z1sO+j+CYpzYXNdH+y9nnpUusFXQkIvNWKAtWdYUDWf61jxNor/h06uMjTa+knvvw6QTlWKjio21
u274/6nUZRXWbJ5qFdzMq3Pz4m8ZGIGWG+nNVJg8adVIVv6lK2AYsYyuq7GA7096AKWZoAq5kVlC
Obv1LoSF+wvwPH+gE6MWdfYV/MZn0HI/+Fp0f8ZtZqExF5AGmCnrITFpRzFhCcCf/us/V2TUUgRH
pl4v8L+sZWEZn4Yhl8QjcFKGNQ3/TpxdWCacZ+UzM6GfrDQ3YvZep2h9BGV6IK1zJ5ACySPxkq+A
znHB6C5fHyy+KYTcHq91SSvIsSvK9ekd3m0vlI2xjAJVhzdkjHhwFIY/N0nwSKNEhezAZm1her/e
fAamrIgsK/PKs6Wqjgp8W1yRArb+nOtopUntRFIQ5/yI5trBV/IqXn6re1I4cTJDnIbJI7R6P/XL
7TckgH0Rx+hpF1neh3W3C85fiMATfy3aLRGqhREnm+ZV0yRBCw1L67B3SbsfglCTi446KfLNzPN0
cCM+OKjJQtkcXhWeBYsb7bRvjS4HrIHONGo5SFG3ZVS1y7KRpSpDutNtEpeBmbGsfjGE7DDB7/vw
A0CU2VYOpr3FFAJdM5dKnADdjXiVCVtT/Cpa7JokN8GYQxV8O1Wa9PJq0o2LHL+LXq3WZtwrames
excf2soEUaHqhGPNAPk9vlgqj53BRUhmHJmOi8p3Calg/AVhZQeFQtjXrM0LEv5uklnzWmDNCz39
XZULclVvUAyxydSeTU1aeKRumrCCjQEcNfbJ8yoA1IYRkoGiBKBnwLvo5ONRMk77UJMmDuj10HSr
eoWJltexYbKeRS7C7C6owT9LbcjYvZ9OVcvTQc10Kijyi/mVySbCSASiCHcsGh/FNZ4WxXouQm/c
BTRj3AHLIFG1B9G2P/IVpW1L9S/62xd94AZ8ZqxeOYRreZvCHR6b7jkVvjbISoWJwFC4lSjupnCY
KpaKk/H03NFMlTu5q7DmVq/nLrEvNjIu7vx41QZlKRisDoDl/BYQm9wTnkUqyJbBcX7/p4sQp1bm
Q8yaW6uKVk5+0zxSc7L3JbLeEoUEe99LYsCTiTHjw3ShaS6AiRUlb7uCblkdHttiyncvnJ65AvIf
FmXXUn0c7MyfYklTo9TaGHJJ1u1w9Fyu9LPq4rGWRYOeDMwZVd0c5XjL6ADGQR7qUEZ94soQPxlZ
H3BU6doAygbEoIGKSISia0J7g2o54Xzqzbmp+7MEEGyo3c1uFiz3FHJNBDNyAeyljArEzqpgAtFh
UgjEINW5g19hd7LOUd0blXBu2dbJd3OZvxNe0PWq+/yRU8h9nGlVpihXVdR0iEpcRavIzHiOw+by
M0oGAfLx2B43uYi8uKFEKKklMQsvKcuLvab3vpoJ7IfKD3nKwRhdLwgeJY33prB6exyOoObm0eGy
rmmMuqR770aKNAORUztJUP0gaHch8NvOqu8E7QMuC6G1+Ty53wlyqyinRLW2qB5Yp+IqFupydWAA
jOWHB1jmjY87vx3YrWiGgFUsHVKYvTJayI1Of67SeusK8Tq6cbTfL83xtXKBeDBRZQRuhox7fGlV
SjjdnaxcahMQ/17orpzJwM7KylUbGkZZ5NX4QbaNEzw1ZDXRXku8nPPjAVjXPTz8WPvTmAJ9LPZq
C/AW3SMfLvu8CLL1ysjtBiAvCQsx7ZfDCnMcIEvMqQZ2CjkGLn5pJ3/YeJnAmbK5X/K6C+dP7zfI
1zOQxaAyKwSKpr0uqG1C8d7w2k5JDoRAynz8iowZkBOVvL1AhYLURGhyLf8L0/uma+4vddvz8+u0
Map/pnj9WiRxOo2A0BaG+ywXZRqJBekjMPAbZJc/X9oYeDNCBcjO6y/QCK6RzDbh48DJSk74bgYc
FbHpgxwimZiNijmf4853Nc9sYps181XlXK8hqiaZJ9jpPnRNXebc4cURNNb32SYqQxAvqGdKpfP9
bNxZ2q2Q5+g2kT+J2Movx4r5QvkHstro8cUKoscmZ7TQqwSKCSQ667r70J3r9SKHpkghIGivNhe3
DOWfiFkAsjZ6YYTTpzq4Kvu78ya1gvuIGPy7/IDNrDkkZese2t/UnbnJUFVr0tWQTIAmABb2PkSH
PmzAbL0n9csXNITzmhgpQEZ4HornOoamrSyUB9mHsF+FRAAxMFq9GjiXR1dCfa52eAPRuC5jy4SP
5bLlAtBW4pPNMjT49AbdKdBuBtwQlx98eXqH1l2e8g2q1NJng2duvfJiejk8pnhi+jFviixnfAMY
NNzTFRU/aU1QXKb5BQdVLc3oUIeak+2YfBj6NTwxknZAxmv335T/D1CQFjsp1vQp08GXCUuc7FGr
GOCdu77Mdpiy0/z2iMIuWPYsOYfjTG24QOSjPKZZdZEX8SPbTRGCkZQS10Ne+CArxhsCydPAgHCc
k5qlZ0W5WgBhLJwflc43xTcXZw3uUb6wnWUIQoWigooBDPRsj3drVMwjSi82bgGN74ec3wHvzNl6
k+WzOiFS0ctJyIjIL61hGHrYViPS7wi+/oEf9PovbrX1Ox9AHxhBesofSQ4GQxMNbKN6Pc2xHiFE
9SUHnXQcXyVHT/Wgry3OwhlLIxFmkSN0j+EIoOrlTzkPqs8CuzosnYL02gltU+sCL4i52T9RiAI2
WyW3UUJdqAC55LztL+muFJz4J/MtKtb1ONTT6uzxVAJipeeSy6ttRfDw/B1t2WFhZAW9kCozfJC2
32qJCAMYSZO7xNXmikECuQVDQ9xjQcsBNUcNzBw5v1unQFPkZwYvTAaW3Fco2Dk9qPQYQlA6X3Sf
ELIZa6B4tAdKMXvlU/fe4z0NP54AKkjEzfFHupRT0bUbbQmKzS9bSZ8pNLE2peYafB6ChgG5yyRK
VmyBw0De682ZDK65ZFi8ttSIlYXtlD0tYGa72GJ3d076CiXPpi6g4e0t28g369jK7CyRKyuez/B/
k+074E3Zps+YHrc08S6+7YcIqtca3zx79iwZvIv67zFTTJCsSw+U+gv5dLtJZbyEfa4irX5tfegn
EdiXDvyMuRIFvragFF0I5YMKFpzSTIAEswBIh26Y2+EW2nEgv+CHSbYSwvdqVa3+kZDSaCzo2bN4
LBub1qxtXwCjF6lkjDXL8yzsNbCI7OY1U1nFLZQRPg3Poa45x9pOXuyUsK0KMMYzOjfxQmBPf9GG
FswZZLmJfRRYampEyBmPu2hZWbkud30fAwV76SHubaLJPzFWn2RG2OvU02yv6EOQg0WQhTPMow/t
VO6jlQfpMARSxDSi3q/CMiwkoAmfit6QWfGMoPWZCz93JCiXW+BBVGnkkBaaMhGVYmFutopISS3J
CJ+ZUlrmm8M70vah/ydgKjqlGoNhdivZaQp8q8Rg04uhKTTCdF0kzIqQUzKOBavjpcfDpDjBY8EN
A+0RpCb1z1CSQdPhiAx7MKtn4M0e9jAyKC7MuyiLA/GbvISNDSI343oIt7T8a0f9uSaSylzdIm8l
mDsBn47yZH5TgDOppV0j45GSKSNwe1fgyRNjC9Mi4U15xWW5ZhbmBuzjarsxh/yIskL5iDokvpOl
unHHtuMuO6ny3M2F3VUKhVMERFrX88FdKCnw+bFEW8682BQ+7JBJYZdBrLqdS6IcY5VBeTRFuPtA
6KvcuX+23NY8ZzkWFNEe+hRwEfZAjO4XT0Iuus7KbUsk7i2VUj2c5Cw+iNhZJfY2337g29SESd+W
P/WcJMYNTmm5FZhxDmMG8ynWXJylSAxhQHdfpBHNsVDx2lcPYSrA6d6xI85C2W2M4AeLRprBNrTr
fUnqgXL0GoaKzNjl0c5lG8NVtOoPqHsoktj2TxZSSaYfYpiMCePwkWzoBCxLLvGPaoKNhO9x0VPr
OFU8sYhJRzHpoyITtNcr33fAbPchuvroPSBPnQXU+9EAr8itlElyzvNepObLaBxfYCD00SPvwYED
Pdq6ma9rslNJ8DaQEEBpunc30u3fQgC5EgVazBQsXREHxgOOfQYAWU16BoExw0rDbFF4CbehWKGy
LZFqVF6WSdpbY7optrMbJMPR0mHRcB04CE9734MrQZl+3ENUqI0i3go/f0vBkYQ2Rj5MjniIg4yp
g0kI1MbIjZhKcetPxg6bSTi4uBireT685djCeIIBJYjGVvGSJLcA9a8dUao/YKTh07Pg/5GYdj7s
nVyBhBBLPmgFViMmnPNmrkCH2u37F89PLn/wqQxg7GzI9PHkTBPbLa2eVdYSutuSikKvY7jEav0G
+KB3s0JskUdZ5d2NIZYJ+Nmmtfo1iQFR6KKIiNHzChmT5HjfMbwaV2IIQLq8hpQtus12Mm+1qzdw
v8NMj/c678qc2QwuE51VkL4oz6XAQP+BfmMHfNn+LfBbsU4hNWPRCqeW9yVhr9ZFlTJnDfwu8U1U
ZixzYApd2IcB43mhC3yvjF9I15x9+IyyFbXymGQ8DuC4GIVbewPlpPjfKSSOZUWQ0apI2nDZz/tm
nBqTxg5gKdGj8hWpZAbMGFZ04slGSYPAIG+Tk2xe5WEF39kR3BaIKfaZRwE62JYUfNxdy8iXGdbg
OzoAMQwEXW/zXol0hYREDhn4pw4pqRgIUjpTQJd0eHNiIhzK/dDB9wMgIIwc8Z+LSEgbRs0Y3DEC
h6nZQYTi0Xo0ROAxr8YcHn4owu/wBoXoUONR8/qwCoc7jGls+osuIi5GcSslU0mEjGj1vWVSKcB+
2bB+XnuG2bcsojEGxl+QilF4l8VfGB2TpYYG2pSEcW+vX1jfTzlY58WGz8G/vmvI/3tgkMWUept0
7rV4iF036kX0JujVuSSHdiUwWmAcHsIFiWKhwIPQ1YCrz+5DKXHhTNub1J3YEzOgTzEK8HVHvmSk
gR+30FFnl2gEVjARHCdkFGEnzUaflZczOkYnLh6U8J0oAnivf3wyXX7LDD/42dWQlXR0OHdtW10m
mm2s5O0ZMz+TAGOTaB+SvqFKlKMaliT6AdP+XOUrw64MtCfH8w3M9c3MzfQxd9bL/nSBTfBAZlaq
AAB1d5G2fJB/m/JTOTILGkFmJYA5DHVmb+/JyjdXLIN6Qj31uTxbgX3fFsOBE/hZs05Ad7SkSNvr
WNrFNq3aKJB2AAdNtg/O95p6OIfyk8Nko6YrXs4Gp8ibPEu+PxT4vrEIImhvUVoT8jgVhNLSHiq2
qs10NOP4MkoZgdCGAcXAiMVLbSMPQ/4mfPZ6xg70yFs05hVl8GMhBZ4kpXK5JZDYQN0BbyYaPtw+
uu8/P1Ngow38vQx7BCYOVVCshe3UPpkfWacgvz9a7Nk5L7w/S7ijGp5Tw+TzjN45TqlsuytxBj6I
C4OhUCX3JMu7U8MzewN32GN+KNISVxXRudnAINp3p1twTg5id2h4kVZfw4MIwR8vmXv1myanhrJe
vOJ+tRX64kCXVMUPa1Rv8KwVmub4IF1FOWhp0pueJwAcoXSgrj7aLBk4n0NPpLEJCmH4tXLilLBI
uS66AXFOxiDAgLl5Bb+/BJ8Mjiz7go2pXzmSJoAAKvdSOaSGdPLzitCkeclZBTJdpFjUDwPtnpiM
p/VjL3RfBsERd2FB1IB40j2ihOSkE6Cfe9NI4HUR/uA5fi3lrKuF8QFbxJeT1MLzOj/UB/oAkBaT
uJPgEHpqlMewEwAqZ4QZDw45jwbZ+ghW+DsKF6JTJQFc3t/NhPPeSBSAFLcBpF9Qac6rrWXjDLW5
ZWJi9W560Uq11GKuW/KA9zGerBJAsT65KnZdUgic+bl6ymG8doPojdqG4qz8TFD79YoEO5EMWkXp
qX8qZwalahUQ7YwFH7Id0vYLxyLopgSFMhlteXT1qtT7c+Dv8N5z83HF0KdPEKA4nTWMhvmzcaIP
D/eMkmKMfI/Wr8FpH9iqxla44VrVtScO/h/ha9fxQjZaQnvzSInfwR0/0VbzfwmYmhchCfT8fhMY
PFrl26fquF5J6zxzZNyr8iPRhMAkA1tEPh8bHGNMmShfQPx6f4vAeRy9WDaQI8NbLW/pLBqDFy9j
f7bTdP7r/WYwBipDqEzjXR8fbjqGZYhq8dYlk2L9janPPR7nE6cJvTTofbYjlH8MAgNn/UFgPnFN
Ub0rRP+RvwLRKP1gjMPQFA0xvllEI+gXH+yl1T8U8xwotCjRn0awrBMbd74MEeAa5KXmMpCDvpFX
fVFDeNwvuCmKaLVTgRTaT/4VhmJOQ0d5CPvRMyPZfCK/pM7w3ZP/ls0235FqNAptt8qf1bimS60a
cbxJlQ+oNfQxUWqNNJhEz6QisZnJQoExfEJUGG6BJlzrHXbByZDbtpWkIcIkGs61XPcVKLGhbchv
5sbx6/4yFk3d8ieLuDNInBiW6a5EBIt00N/a6oyzHhkNWczLRYYOofNuc+ACu+Do4MWUxN50uc73
rd3CXtw/ZI0C/SSd4TjWGoxRF6ydM8VPIXPknhwLGWDaWkD0BKasDr5qFiqx7p9RUNtJJIG3/1ZZ
ggixhFLsX8HRUoURBPANVFdiQC8r5GqlmGdjuJ1F24hQl1iUJIjKX8PuhTQJ7TCCSbiAd/FWCfEX
iOXxGRBNLSmelPCKRkopiYvd4TrdMj21eqCSCJhE/9iAZooOf9W0hH3AevJvZ8AYXInVjWnz46LV
o6jmWP0ieRF/e821TD7wfyfKZEoOHl7WT8gWl5xUNU1ubB66RNlbtT5gOjuzqOJoQn/iDKTJxn6z
1JLoubHn6M7CIds+1ympALhBZf/q57wRUuUBq/PWqcg6n6ww7qBPWnaY01ytPWQi1562s+C2jBNk
xQTsLn8nBw5HCy90PR2jmlUJIS0Fya6SU9WEAPo8CWdZepHuZ+P+9P4QCyAqicSUkTZA4r0WxS5b
SABv/LZfxvSQTx8F53L/L3qfsh7oaaCt+xpZsnLpHll9+XC1DkDtDzuIurLwPJXOxPEZCQztSsGh
EtnBHDYYVwhe5F2q20v3DQEKjx5t5ySZVWarGcm+G16YHemDE3lLJxxUlHDDe5PQFKCG29EV8sX6
GTcAyL5qSpwDVKFn0hmwxZUJxuoX8qMhk3wibGNxpvPLil51+mbNFivYx7ozCYEuQf2yMLHK9kVn
zHkOgs0gju+zd0MqxXMZHXmsPVbkCfPdpMKtzX5hnZw3gXwFiuUJUOe0ikGbQzkolMfxWEdqWuVf
N/nBkDDesOk+xLxwNAD+6bFO2IBG/FxTxpWWdOToB3dXoN6OnH+mxHEM86IjGQHpY/jezNhVljAi
xeF55B/1m7exOxHc4D49McEcxaiHVnOKBXuZ7Ht3Upvi44gcf3hDkDlo4z/jz+mLkbbPCS0g4mw7
kKPnNwJgUZJaslAgPPqZFqhzk6tJlVWKuBoqSqD1O2tjDAhwFYeUr/SCMLJJ92TOGCUlZnhZD+Wc
e3MsyCCGTsg4P3CwoBuVfeIJzdkbuez41HEqBbibubJVvLmmWeiAqb5eNT/epLTJ7MXbyFdjqOCV
qnD67jL23ZKMyNcWVL1tyPvE48tbrp7Hvm34s07Y+NHbqz0FSjrnKn0lMjQy9gq9VD1z18uQbpDG
JdCdDiFCAJ/KQmUZ52PgG6JrKYDhwd6PVy9LU6w4xWgtaA0CwjoxmzNOgKokKes78ojuex23BSbb
xGPdef2W/YcpYTbL8NXJ4aV+pW4Le1BP+dGw74eRrwAe9c7fB0TpaYd6gYTQn9GiIfUjsFuBmnmC
ntqx7jOFZvecWTRyYywmLQ0TedT1FCok6/ckp2XgmBJ82kNg26t2olvA4p6KSHAT6ofH3RJH+3MD
WygiVoPCmCsu8I/aErT28Pwo9j7qvDfUZTSNUkF1BAVFXR0EHgpfCVS7xyJczDxuaYNUWwjKg0pO
BqZ9dLzxdpvIJ8+b96BZHoY6ejnskVdfeIlpd04FgN5yIlRf3kqtJbozs5cdyhlWu8XIhezeR9e+
FSJLKkqpKBTjytcLQ9N2oe2BL/stMpyesjPlS6rL8iLe0sJr6l6OZFcbcPicVdV1i42ayBZqTZO1
YVxXhNW4NPKNTFXn9HJpMWhBw2B/Eq2Zq4vi53yEk++LFIeB3Y7hG1YsY3YjnXNGqF2do8ZcR9r8
q3WKJhnQtHIFX8Oj2oX700v+H//8u9+J/y50mc5qJyuzQvGe6D4zMr/D1MF1EiusoAcl+I9Du/Hm
AKFIdKn7YPbuyRfu+Qc2IDKoiYeYSO4Sg7+R7O6WYy2KaXpVlAHlMCZSC32V1cz91AkX+6WH4UCw
jgmNI0MOkBaAlJvY802f9KZLHQvfi2OQhAvM+7hEY62QwkWkYM162UmGpRaApSH5mqvsh6U4YVb/
O+0of7i8gXQksdXnBe/C+825llLuF5sOxjYBVEVCXYacW3LnEQHyLDQd0aBbcE+81OLBg8LJ7VP4
wDhNTNKTAmzALLadl1z9riCBj/cKjVuHiX8xfIkRaRM9DVhsScbAUlYvIWOpBQMtiUtI7SxoJwIJ
+s1rGcqo8Y5swFS3lbfMtvsHwv9BrYxgr9Qa2SpgDCzpGLyYIUxxvl0oHkGgO3HfxyJcjklExAjV
ABI1LBH7F/9PiDXW19DaMBronu4oJydttzKA5THFhUjXiSRE9zOB5OvNZBWg455E4ki8vll0ycgr
Bit5IOmbEb6S/Mb2xlxSsi7TmPzjkJGfFEQSyAhx3mmlI/HX4lyagRkUha0qxSaYuT5b4BLO1c5R
Fi0RWhNexZ+iMqk6mbMQlgZH5GbFqoJg1sPA8yHShk3tIqn+NUHuXXpaOwbIDcYBI7ph4A/ep96x
ngxQXySUGx9+jpO7tGXKFjPF1ohQqlYtHXcLoiKeHYL9TJiOEZrtwRImRxakCRSKathCBvhuhd+f
We/3IoNwwrxegek9TohKUGrKvLY+71bBB51ILPyUqSBxCRNSmZSL8NPIzMZxVxX6rIj0CIUaHqDn
DP+u1EW0bPnv2ddRIPuv8JyRo4AEwXE1ckMPHPT5xGNCiJKNjC06fAQkYXie2WsvRNp2xh2yUnP6
Otiq6zePQUYfJUxZNyp/gzghC2MJhDQFmAtxeFG0o7XCpaph0RWxF8jcHf+ErlY80/RaW5jjKDMu
chPJcN5IS6mfFI32n1NC1tfyhazZdjDDvwCKypZTfhEDetOW2Pqqf7h9lSqI95wAuQBh/gsSjEMX
2vG7vYsfWXqReFCvdUk/ntqlyyySD6f0tYXMj5w8ny3k6QmUZZht8e9OY7/bPTJKea2jC/adxpYt
M1p5IHnnGZ3fzYorDHkrkJPMskJkt2Y2t/CT8LZbiQaeMkOqSnJz+NP89szAbevwhRmWTYVKJIBS
uHvjEjzvLc3gEkIfDbRQX4v40r3sXMNHZzqS+iwi3gH+f49YOhNJdCaoiYPDjyJjDMc1TrKgPVaS
a8hF7+WtFuQ9uqul/imfKLmtrqOV79hTJc3uN5lZp236BOZMgb7zVi5nfyaCT8RCODGqZZ1EDsIQ
nnJ/W6/MAGyaio3RB+w6okSsOgDX/bGrcAnQP9nwkPFDDTiLDkzWRdu9nQHQ7YHqfKoztnHELYca
Psor984jyyIoBaQBAjkQNuUEI4Eq2Atn+Q4GClwoeFv+KsOX+CYnsvfYqaEdwYxrNK+uNRdVBZ7/
rCLrG8/OhhLL/kdJY2IVc6cS/ZUvLK+7PTetnmVGTRZp4s2GbJmiuaUInk/+/iV0aSgPmZw+ICeV
p1utvO2qRAF95WCPzWhFtEA6LMX+qu2YilyoHwVDkETLfJIDsblOojfrfJ/Is13OBmV7/YYCGOOm
Af5uMlvrC/aqIyBgN9NqGCeE9auHgz8uvSTUZMTLPBlHqGlUxJNAa6u8s+5YuEb0zbIqjT3FgXY5
zM6teztgm0WbHirjoHsW5v3K1NbxVHNT4OcgQoXT2xv2wNytTkqzu1UbFEkWxA6shP50FJ+uu63o
Pbo4Zf1TGHbtvXEEop7ZwujqcM579xEWm5kV0HW9f448JUKlMH1s+LDHdqyWk2pq+YAEbZW7a/qP
loiFfCrgGDvak+8yonpfJ1hZ8X85JiXIdiQpLtLUJ1kn0MpNcAYKcz7lwJPikJVjWMuRefv/FsLS
KLyQjoaM+3np3J2583hYZRDZgfBlqvllgPb9FGZz7+jxwl0I+rbYfAPUjrYinNMnDC8RQHFBKg7k
uO+A+7Y29li2Z3Kiowl6z05rupe4303dZjF/AyLStj1bj6BeGpBaOOYX1fALtFFRsJhhiRLEd9r3
oew49r9VlHtw4wPW9+WOXDrvd3IyUrzsjH2q9LWDmS+BIhd5yv3WnSavBWo3ZTRpuqGHZPVxrQ9L
b9gQrDDKuC5d4sIyoAyAu25uA88/d1hZVkg8hiN1rw+gmMEjWxo4L+BDgYj/SXMIwm7sUDF+n7Lh
8AAqIF9G4n2JyKIGRjGcMiAKNEKK8TNDDhkpyX+wfXNbnCXcXCLWZLUCav9YoFcvSoVZ88/hGpgs
rtpGawsFu+jWxbUnoxQTS2bm0yBxt0FwJkUX809oKMKWku2yWTh1ZuTkzZ8MuvA4uJ+YUjBBobpb
79l0633lP2b6h/Uj94XkrvN3t8oXIblPmGp+b+T9FTAQUcSeOjdKOhGWUqR2SgxEWCzEu0UfWoGD
Z8Nm+uzL0sQY1nc8xvYolsrhvfHnc0zAGcUfEBR2wMp4aRNEbyWmIZQRW6s5710VDXprs0bds281
ie8K0eynApmwxR12plvEaS+/psw6nD1UAOThQ6curr1m6Y4FCDiYl5yYRjqxrAGOJ1AS4CX+Q4D0
XItLXd/7OoR6x0HdoKgCtDDs6I/WesYOB7DbjcpcXv3jlSp/c2Q582dVRvGtlNqvmD4kt3WsF5DZ
zBdV6DocpjAcniTWHjmVgl0wkAv8jpghc/Qwlg1ZM/KUdSgYBDnutzNGSAl7SJLL5k8x1EkkzCcf
zZcR0/gMcq1zPcIf7rBXqi3PAgbSXjhBxe1c8sD3SVdPV/ql24jNpo0G0Ls6DSNNe08BJ5BSL6s2
aL++CeyzNyP6RdRCqAnUZVgCSwQJ8VB5OCYccayqj9DbuSS9ty3r+hRgEtvifSgT1yMDuihc6aef
VlUHVhCav/KvU4Ox3XgEo2z8WJ+KtLy+PLjlz/iBxEiHehRR26NTI6KnLrB6GHZVWp6OZ0486YTb
f2jPPNOnvZbTrOw60zIln/+knvyNwbHU3599SqUcArc431QS0gFhQaevgPd53RFIOweLBrOD7E/I
N3trFL1hcVBk53Q6X+6ohDL0CYrxGky745gsDGQHJE2c91qfXv/HFm/VEw0ZrYI/8ogaaOnLPAYZ
/AwqxdUUdBGVxdyA4Hkg7UZOadSIBL22XZSqKUU1dVlbJ57maBsxXK9jY3waJFwD8AZkDzfqWz1I
AduGtaV5Igw/nWaS+BDnTJDYy/bl+VGWMpbTpSkXRZoNtOCqQDTt9vfYLSITTKBVqOKVy7AAMhYy
l9CMaueJ+IWRZgMD1ava48LJZUuR6pL3AnhW214xWuvSKZ+S3ukUVTAimhL+Zbs9hEfK48ahhoKR
mPMcW+J5K4/3Zq+MRFAH5ySVR5owbAXiveK6aVzCz1aaS5PRh142spADBqguPm41LQegW+cIcFQX
f1GReF4dLMaHDcx7j8hFK7OUaS/BwgE+6OcPvl0maaCSmq1xiGRCmGZxT0nZ84AWl4ojQDuk5GCa
MMPjWODWiEkXQ80lOgXuqPfjC4VcRylaVdbE0zi4+Lw/XfDTzs0kk+a3qLzGduwGk+BtmyEIVSwu
86dw8HYVAWgNxMKkejYaYPh8DCdwYUbwspfGHJsRz9m+RTeaxJPMTTa41GuvCWBvN8+YssOph992
y9L3xw/WtIsPWV0XNVcaqRdlAeB/Hk93DzAA4aG+e6UD+Eh7XYGR2yX8Opi9bMR/uXM0BvgqiPyE
AViTPzNKMBzUDqr/g2S/oeSSMo6Hd6gWq1Iz6i8D6Hy4ZXnInx3CoZHJD52QyGqTP3tZtpIryzKl
0YQdoPW8CRV0a0MThTN/rnCR9eBTzhqFcbxXp0iyCCJAIsm+iDph15icwJNlq6RTSQCBKzqo3ZJ4
YlG4P9YTS+dqx12McGvF1zaUJhQGIF4llr7b2oPbh2iOKjXuoIsftDOMDpMAQThwXjRNWtLiV0b1
zNRd/xHbRrHmVCyWd2GOi/jWFHq9THdxxbu0DPZQVckKIfode4P4wnPT/wwLbpPnwHWauFos5xA9
+jcIvKeLdxH5ZMdx1Oa+fbV0xgsJjMS9xI5ubnQJdWWJ5LFQ3nF/tyqD0I1mk7jLV+HPVCQX7UQf
SfzTqpf9LsDRxqdDyNihXiwpt9jhumytmjQCnuZO5Q2BQ1qWiJ0N+xwbTpVXrQssxigO7cxqTg1v
HyT3Ej+ePYppkXG2TD+xu6N2A5pUIvpLD69gPqyNV5y4E9ye0n1rgPW86HqZOHBYjl3OVYrBqSdu
+4yKV+NfAY4QqvLiWc2jMqCEauW2zkHkYVFA7LMbjENu76NWDVk5YEUsOF7mKq4K5Ji6B1USDua5
Tudt20s/4zYeSXcHoVOD96NnnAQea2rLsYquAA687dRj4mBDGe35iqnpiLcPUsWBUn8PIlkjfIIP
crm7i85HS9txQ8CvhdnRvMX46qm43QEVbX+XBiwE50kO1vqjjcn0n/3fNsa+nPhh4ipQkPSz/ylm
cPV0tLzzPqCbsAc/S54Q9Og87EVesZVD/I7x8C6M6xVST8raIOYPBRvUPODsofAkUzCAomVGJKzY
ZmMZJjLyNvpWRHgm3IOB3W4OMzNXc40Wl2g+Orv9zxQ9J4JwIuJjZfFcSj6ymt3JnmQA7d3lRh68
0tKow2H+XPIgl4OCDX1Oij3n4pqY3ihbj8DLD0rURQp14lk5cIl4lC+UCRe10NlO/Q7JPkwxiEP2
mCXA+kKxsKHzUeEsJFpw9MlvwS9RX8WiIRzAdYxgm0kI24h5HE1UCxJJY8nIgcdrHi0n8cNJuaWY
pyxaB28LZk2ld3wLkMpQIZd2YaVlcwZUYJAolPtQbtophM3a/ayhwRAfpRcOawnRqpFdbp6AMj2o
qp/FVT9/J/oYSfh+KThcN+twtIla76dVGGuON3M1uucDJkemMcsbDh8BUaopSCXBNWt1KqyYAJl4
dWrepf1IBa/9/xPMcmCeI2qJhlA3RIQyq3SaMeqTQUWL7fgghnGSInEVNCHeI7yOs8IVcs7kAU/M
l6H4/suAN7JmW/2u8neqau/WZXzZTtRLyM6bff0oaq/FxOf0/4MG+6It+UpmpgDtzxsX7HJsRI+c
SLKfzlTQ/2dEKB6aUnxG+Y8HFz5hknqCQWH7G+pOnZkzWtfxSsL4/qI9Fo2ldMykhhZtfVLbPKQG
KJ8OL/qy6PY4gUISQpFfGLCOzFff+Y8rCmEFUnYCOk6liMo1LzTJc1qcDjIY7V5ni0D2hpkp0pQQ
rOpSAQrRFKdxrfjk9e4MnJVf6EiO7AW/59ExsucxDB+lwzdz0gsBvFg83T1FXvPuyBKDc1VtcNA+
o/gXGeNJo7167YpNHK0rgiBpNzJXwhtNTee2WSn+Sq+VsXxIlWsIvK66Eh2lOqqLICNDcEsTCnlw
cABztFxe+AiD6nQc6AMbYTdffXEhYSfhg6kGCTWg1euFXLctZjlwkQdHStMAWO28z4umjGR6Het0
1DhKlYIjkLpdJnWL7qeeyCyks0U6omzMTTVPXJxqHzEasYh4M4zjgAw+hhaUuHKP1zGNIEgGzUG4
Wkzo1+hrbP//Dytrlg6gKQDq6WERYl9WHI5DuG99fKG7ubXjQ+jWilM2N4XaLtzcBk0oTutrsAly
Lhx33uT7WJdtvwuyqNCSpB0WnofMXLsSdSxUp2QPH85Op6DSZivIBklqNKFZ2iBP7vSFEX0m5b4B
6HOHO6xiQh7UHMj8LfwWoT1iMQVGR9kF5zumuHyZ9D5dZPuWc5f21hZGvs1O+7fR8IOY9JVHop2D
6ZaAtnKPyQEq4kTynHflQ/okzXFdVGGSA8g+NyUrqso49uLpILPiNazbL6lAA6JQ3rqInXp8uDTk
qGVo493n0BgMD4QRPOGdRhh4Sn74nr7hkW7GctbsM6nLWjIflZdCR7bxtZ883jiZ3FxQwH6k3/n1
5k+oaZrERvB190kBh2JrpXe4Oka8Sp414I0s3fwbatkKy0Q2uTfRtMZc26Kd8evrkz693ZcBcUpd
WUbud+SZrtAuHaN/biRTvIp7ly4wSxDqaJFT8is9a9b+WIy2w/e0T7EgoXTu4yrtoG5zQ1abz6uz
s5fvP2I96V/QcJz+fIgIJwrFzYjz+UbIDQdLpt0yF54B0VpCLW3DjMZxsrJszVJMU7oWV2uaiyfU
e7AkGZiorKud6lGm3ZMhO8loBqWYbtbVvD2jzCokLokBUfJYXioiw/5vIdRxYh7UlTdmN5R79DuP
oGNACmnZL23kbLzhinBUhv+fe4alJJgYk4cGcuwAb+nEjN126iFYbMkTIyrDU1Kkc+taXhVwZK2K
xly2p9RLNbNfWIH2Ld/fJQVIhZ9zCm8sjIHlfTdWV6UtgoFhgGj26YLS/MGW5Pws3fJeoA5XR/WU
TqQ74kX7wOCMeHK+meHL/7q4qClOjToWhPcaM2Fnh8DS707ftW+D06JFK1A67TPbJ9W76eNdaqIW
agBdnHNkT6H0rZsU51MpaJYWjRq9WBgcRS998is60JkkRu+BvZ61umSKv8uz9wJDmvDUTZhNkWjl
KwWwB4pcJs4+kqgVQbDPX8nyC2q9BWedDJ2CkqwTRSnsbyTlQUaPg3dbjMW560ZF+pYsdG9+UL2l
NA6R1RYqjNsKRj71pUg750CCCA0ruo5qva2b85lfy+rVyC5b908TJZTBFlnFzXFjKUA6U7hsMbN5
zU0Q68kpiAOve8rwAAOkz4GCHon2W8/vK/7zb16RURd9nE5A90mENkVveAGfCvrvA9XGCyzUfx1P
KADBrlAMKzXND72+lNRPoQqnkMZA1l7FjYxMG2ykJzbKzTP4Ko9M1P7rIpL7X1kD6ndbNZBIdRW6
B0IFMZmkUkJuGzuJgpUfBvXFGs93QDCuHOeJyyZa0764rYpHoqDHU/841Q1Fwg9iVAjyQMfvv+8g
R50MIFs9l3lq6YREB1cYepUqGrxsdDtbVy9z7GN1+4dBtcrXfzr46iQbLrSzNKAJGxC+cmsG5OtY
JQGgET0oYMlSDMyHBdXdT4AJKz9iUA2omz5ZZUMREVd3WrJuGvTYQgOs92i/YUydjxiF6ECCISMm
5ToB4RS6fOuZgsMFjuJv0MB5Jbvn5E97BlGcWYiEbrG3GIPuSqmkEmqsnwrIzj5flU1Xtora1Ze5
snWL7AaR/lufTfhbjntP9KydYDUrgBAOh6W1HQfTuBmlSxy482jmW33xRp9N0RqNsv/Ox5E9W6jQ
ow4MEf43VksPQHdD6xj/dTkEcbqgKHcX6y377AylCde2myDx6W7yq082YiPU67WGxOYlq7KdFF2Z
Fau8icRsdElBZOWWpun+/FfzhFMDefRXoZvR2ymCxd9TOBrwbhrsf7TrPoypys9jWiiSR1CnzrkR
EZiXm380tFc0NsWFc0lJFEDfo/K/5owIkGE1gZgHpwcIyY/leYncyNBWzTo/Z7oncIvzMoM5c3s+
GtwkfafwYKgWu0tif4TzIogzi+1i3Low2bmCzkn2bFb9D+0qmLO5u8/ppX6C8uz66JYixcqr4x/X
YBm+fYVPZn4mTFLOkt1LgqCGgKQSvKDQFOQ3wfb3FrSF8fagAcMlDOxCIKMs1DJYFEQ2wDdTaGLs
GZ4QcD8zySfHVRrLrnICqNpnH546iE+DvjRhRTNBX1rzjTr8060+u2UwTL9FUj5CHs8SkqgxJp48
1Ta2tAxNZN9RMLSKj/1NAzT5Ah0QVjwxay3vkmkALv5wAlEO7XoZ7VN25w/3Ho2+QZ2y0Rq55DNJ
fKWcae6QMVdzJiXeV64Fyr7Rc8OHdGynDU29opNxnbIbHz7LDZRe+9TEihNm+OQ64gOeKiHisgCI
TM8OI5H1Wp3RfU23MW1LPl8PBlKQd/YP+QIB3uDMxHMKHAe+OWGmTA8Ets0YHpGWftioadkMiDU6
u84qu2w/36uOBNr4/yh4wQ8OmdrqJd/1cGm1UG5kQoPykepjDdl4uxXkrA/8rxXOB1bbyDCj8nqZ
n4pWpBRtjjFyYXotRchuxvoOMNtBnMRhifsxG0XdnkBWH6aVuU6dkGZ/MVwZVAFGR95efD+QPItv
BtuR0d4WYHmnkURdHYYj0eerPZwfvW2OczOUcxLsB+IR3hTnnX6zA7HrNHdMBZ8ssshlA7zKx17f
kiPBRgF0oToMCDMSc6ae9hRUK4S7FD+Uf1JF8VMpVWclLP+ZMSDtujI6T8sIcMyHSoklbleO5PCV
n5Sz2RHKHG2S94d2MXraz66KLDF1leDvRmYXtd05hMLRNeq8ormeja5FwQwGp5kWdt0jFsG4bI0i
7CZr++B7yicsPnFk/O/rta9k2BPn9iUFBnbSB+ac9DsOkrCg8VCBjXYwrmctA0PD7N6gz2xTAcx3
mEKW9bY2B/y8OhbeJogJb47tLVXgYqSiGQTwpfTx82UdTYP3Li4CwUVGo/bdbv90La964LEyzmkR
BK1gY6Lg1jqFcS8OMfgEWzEbQGvV+xHgh8JSfNnEhs/QtkyIoR04gak92Ohm9DwC4M29yH4JhQAE
t8T1H3st9PFsajOV9ya3eLCQg3tYRFyYivr+ZiaxjpHx4GXP3Itu28lZ4TSwdMhKZwpyAYbWh7RK
UcRXcjvEj/EWVk0jSKm6HkqhrriF1Oo59qv6ru/315kY474kEe89gmA95y7hteaOwo8KRsY5cIPw
pWEaZsZwDHjJ093lYHSKJ8MfcFUU9okEBtWhaAS/6x5aFHUceHLR3pC3negUoNGrlQVMgAzDrMc7
+2A7ohvUQNyAA6MNZtsvZklJf23mykflgY0DLMhiuxqsNG9iIk+nempow7zrLQHmyTfE7QuwEOAL
YivoTES4ZDpWhR3Yy5em/xbLw9iE62rEa2S7rT6Y3nrgFzLNqYPsttjv2HbtXgBG/KLsouyHSc6k
xqtN3pCQXg1qqZqw/PGo0VDAnuikBwqfWpki4+bCjcHTPbtIfn+/+jlMUDCE2XO8F/qN998XuPgw
+GmLkA3mHev8bd7Ui0y050oKbWhPvIBBjow8SQZQn1KckMD9Ttg56tYoQwSm5RResiiVVQLq5D+9
c6zAhukRxKK3VYE0CmaaZaV2mtM65ZAha2oLAlEgtwFoAsrGb6K06zI1W4PaK7qbw0dVTIfbuvRX
UN7+yrlqdkaLr1XKIB/qRY9o3PWyf2SG0q4uhZqBJjIrVLMPYxobYv2YJ0s+sk7h4oxTU7LpSn6i
Vkj6QajiprQ7BS/wxSTUA9VelVgE0+EZ6frFTrAhjfV5UwDMVC2OS7rW2W7OD5JPeXEpyQ0LacAg
M+hy728wCFfCmabpQH6vPW/B9Dkm83cFy9jh4zM/jalilZzZDKM79IaBNTZfiae2n9JBY1OeHVn8
DsUOrr5Y3S+vGv2uucmoww68G/AdJFREMFCWqACP0TYqwEKRzJXK+K6w5FS+3TW+V04BwMIlll78
VggROhEtGQLRj2ElNQyQ6NPS5MT2P/aIWCUmnThIRupgEDpdRNh4g8d92dPW5KQX7i2ye/jg/K7o
osmg2BgdS8FV/l8JRie9NEQYgs43GAmkZPeKyj8glfKHg37+jrCHwLi5l2QXSzJSR+/+dDSK7UYC
t5N2nXpT4dMHFJ/jYHL+g8yVkXU6A0NnR7EBCAEMzLFcBXsn8/LeHdfLbOHvIDXL4otNXnMJnvuZ
MPMLeb2A5S5EJCuxiwbItWISjc0Yo7uIz85g1cc1cTw1gG96AKjJuZ2e6VbIV/mo8oZdI2muM0hR
Yg1gUHCyUKVxlyWYQ3uCZCszmlycUdC+Aho2rBxdl79UB+hgSfyK0X8RoDGkKaAJRW6OYnJSrLAw
vtqJG4JZM2BqfQS6BgZvh8dyiI+fpSKEAAPILdPrB1LcNgMW0keFMlfB/spH27efo5HeWJkvQWu5
25to6Uwqz9e+Zk7g0LxNjpv/79h3jpO0ol7csA339poyWGKJ8BGfN1a1ykHIImAERKbWyMx49cT8
pax2+CaacTodgz0ZaylgAhCbPrJozXvMm7hYpLxTzkM3RQpWgnekLWrqk/5Ne/U05loR2vyQzGlD
KgObvVtMLUYLbLyxAjC1Urrndx7o9GmlKbe35QlG3fPVtobzkBJYi9Xaw0iwhi6xp2RhYYUoh6LI
OwhinAHEmBM6A/aJz2eVNWSbdBMAexTsC2qwscGZIe5b834Z2VGFrT1Uqt0X7yDqAw/Vtm+YKFFT
T4StXJRTux3u467VI5zN8f6e2BSxRDspPjaKsKqq7cm3mlVE4anxkXzKF4e7YCNBWi7qRqsUd+lQ
1BSRNaXHoho29Mtdxrj2WIEe2bjzDn8jYK3gwAE/Da+hyBa6dDfDYJoE/fcfRCB/+FuSKjU8p3DM
nucw9f42K2nyhcxbZSB/dspZMgtkXNjPCrNbchJ3Zm4+PHzEUz/me8Le71hkaLXk3x/x4J53eGEB
UveDbTrttLd+Daoa/9Nr+xwrFvk0blAroJ9gKv5HtcJxK3uG8b82f0nomvbmwaxeUf+z6073c4Ji
w31UbtYlt9SNkEIK3N9U0PpOvOzPIbU2GEVf+RZy0A9Wgdl+lZnOW04r6xfNcPH39OfDhlzdVm+S
KW4BoARt00T6+XN5v0jRmHQCaPdq8Furjgqlzz+fetW9iZgfkfPmL7zc2vvdAVkAvhWb0K1WumQ1
oN5+vePqHbwQWa91O3rMqof1FbzT0lXYAftzKxeG0Y6JCn3RLS8b0b9hsFRcBFZMBz4Psk1DAMCZ
aRzWMoStonVPJpng7AJj89PQDA8Vl1WLbfuutVbmomssJcz9hXBgsNQm86ijHX9XU0/H6+ZdlLPJ
9cnb7dkMTv/NCsJ8EOIs9DDZbqja9ooWbc3MgsGDADevM+6lMjKaKh8QguCw1+/VJ5a51w5VSL2m
HSG3g+9Mp6G3tuISl9i2VL1Qo9si1du5YE3++xUfnXsuJGdeGWQr7r59KqKmgl1ORGtmxXwjF+j7
Dk3DURP6x5oZoiPTHDefkQWpcw2pkATXQXuQAPx/a/NN376p7IgKa8Svu0eO2wWqg0IAPT4RaUAD
mhEsQFrys31gzwRasrUwBWL8BGAVH/V2kqOvFOnd4ZCATqnvw7EBk3kH7ramKURaYP2/pQjgXiXc
3jeSHkw0oBqQR7iSdYN3FRw81Ay5QTBwW4TrA3Ider9YOVk64KIJZhhomZASzJ5VbF37I0aaNY9e
8YkIoY+2FDQh1Yvc820pdbqyv7UzGJnLZR4HrcVKTM4yWQ0ULAM3kQa+BkuYJGwNckZwRwEqJPuJ
5VkmxmfchgX5lHkP/4LE2rEwni3DOp5r96mEVc5MJNJk1rzwsAtkgVyjXZ+LPtPBo/CONSF55Arn
9TLnGrF+rda9879bLcuumdjlBBgrFAVWAFdpd1l/wXIjEKkpeIgrrU/DjXDa5Z/NtaFpTHlsVpr7
qkEaa8SBgvwMDg8vUWMZ9yox5UowyU4phgS0aMrlGMADvLE1W+BHPOp8EUJiOGgiPtCMKyYGyr+l
ZkXlOO6gw8w3/g7zjRfucFLkaKBBfuXH/U7dBOWDQVDDV1GLUzdLvQkx2PXM9TNnxwkmvHUq0Wv2
A6Q7EygpYDA5a/cFJFUylzFIXod3oqBR1DuPxP7M7i7s3b6bU+7Y6/1tKciRBqQqznIbEA/GxhN4
wFCV/5ExUzk/6/0NCf663CmZ0dpiaEK/RYDd7eYwka7MyYUlzF7HWqfTy+qM+l8a2+sFaHT5JqB9
tt/LBvRQ1zu1TtmUHml2ih0ZRh9ncFG27spHaddSb7ccfyk/5Jr1FnSA99/VneH4Tg3HSpzmyiDw
QigCfTIukwF/axogeHEvSHCeRn86HYS9eQ8orAJ17ZalEPTBs0p4rsZvTMx86cKvCOZE8NtW5PK9
rM1wM2pw49fWEZz7QxeZ+uzF3a94OWvEV1kNAFLjgCG6vK3XfySE5wgoh0zKTmwsvWK6v7FQhyn9
kVtY3Hn1X0kzVnGS65DGtj+bTzJIC6sXOdBtf/9mjpTRjLYeuxeJChwWGMZjm0qCNM0SP4CHg4A2
OepcEiX10i+oxHWb8U4jlt6VphmDJbj21KRthyVdVpc5WCl1EWBRj8R1T0aC2VMTCfXYj9JOwu2E
OeddeK+i4qWsew0EBrC3w/nMqPltqw/TGmkFviTmpVMWyXQj+lRfwJFkGmDkSaePEt6zT/RjWQ6w
SKSHBa+gKl4ZfgnwEyZMn2Jlh1+NNOxEKgyap6la+vICnPG+5c65LAjbVtCfRVLcTmTX+5Izltfd
Q2mF5osPUUw6aOrvXcWl9dGWI7aOgLDpqjQHR5S/xdRFeUnhGx60xepyDTMZj3EieP+Q0i0ot15X
o3KGd7bTBFILL3edYSxjsjPvXmpVucW2owad2a4mUTVVj32BytF7u6u0u5ivzeL+pkiHhXiQ1MnN
E6+Ei6KYfTs3Cdw6EZtEKbeN8jaIwbzkJD9o+ad8uQ7fSXNFsPBlb0XmUHRJGOoDaoSVapyH2EtH
xgGolYrRSyTa+jkWCyMwnn2l+i11SOZkN0ZflBtSlVs+YYgS0T5tP4yQLhEdDJx957CS0h9yzI00
7lF3jDnJTmC1abJw+UE8d4DlDlX2LRRbE7pKEuYb3BAXlvKkDgMm/rr/Dci/xS0mfUD7etEjaiOh
2PGySPjM9Q0NY4nvzmUzDtKq5XkvT/JwOq1ilqTeSEtoJyBZYDf9nJdzR6UBqEDplMTz7I6G0l5r
TXvFMZd839+8DiW/kmhk48OQDyW9MKFDjbgxj+gdKRp8cXPwXNOXCBE1wNNPYmaUTBZQ61uFG2wG
YOFH/DBhEjYUB/v7nKB86DDMpiDcSlLZYp9IdrgroKE/bF0rOju6H6tLQfxz0VWKkAJgHGLcpTxB
ZC15mEeX0Nr0QqfsEyTG9HdxwHjYnscnnzp7HtkPQ3m1MH2GhA0XqPTuvU4HFQ+mwVgFhBc1lpzM
zUJ/XpP0BEfgD43QW4tw95sjTHwD4YGneemXAWBE+aBNvrndwm+Vgvly+Pktm/X+5CQiksl3uraK
SSGOMua/jLggUq7uhRr4QB4GO2teAvalW/8wEGhbOAPSC0T6RVto0ktxjo+ZypTKJAndD8I8z8m0
Iqw69FkfRnE+pDlBAPG3FTlXhMh0NpX4yd2S5GWl4HC5pDbPY+4rd+klp1Yk5sZswk/fCmruYVYN
fZfXaDKxU0lDJLuC+qmIBZZX42zLEDhVF6q6+lXyDn4a9Yf8L/Cp9I3MAGrew+Idx3aNoW8yZnO5
LPURNIi7ZbXKulGFHWJ1AGzqM6PMyN36lOq67iXPUMA0CrokJ5Tm9clDwM4o9UlZUM8tRI4FCWOC
eyrLZwV+om1Hgez6c256bFTEg1OO7imUU8OQ9Iv6CmtPgyp0xc7+eYxlXHkTzfJan5uwzhTs4ssH
wZ90FSww6PjhXs35lDWaJl6AsKlaW1AeQ51uAT4rKwL3qWi2QaORrREbxp8gUb1dXpfHzJyJnmJP
bcQXNT1vmkcn9KXvZP6Bg9hygH589lK/t8XNy5+95GpjCoegPejM5MYpoJlKVHdiiBXZUyjvM6mM
nQIOqA+Z0zyr+jS2yWGGTl+VBmaq2/2LXxgW06NQ6yBNCrl1vfNG86QNhO/68Ca79Fe7e+VJPT5G
I4NN5/hWaVa5cwgVcaGWGR/DfTLIHl8uknbBwQf4lLOYHeM0rBZWoEJtKQZ0pQT0yFIyrer5T85r
1pyhxH7ggKFs2DlgfN44JP9C2WmYKef6vJzaWJp0vo3HykYZeX8nCl/NmydMhFhVYY8aG4RXANAI
CFBmHDdWxvuuAngSSZl+6LoosbY5OqwoAvJaZuc6Kfh5otHv+e3gNsCpV5zM2dbBOY22EDfnIQVh
/CG6Rd/UtPjjLIU2ftFf0xo0EXle+9KSrc+U+dqZAEv/AiEhpUlrYiGhFxnJKrHMw5KfHmn0fFYU
F6KEP3XaX1VkM8n9NK5K7URFN3PN/lII1/sbDdkEMZ+OBLThB4RMqD/cgPP+9GDhmjQXSOdEoiRP
pdS2hfB3tvQjQpwB8J7H3JXHqWoObMiRxJFrpbNQJyRcDXMtPQIF2hQDBg6Sx0elzkAQxHUFphwu
G1lZ3ao1QlNsVQTYv7lEdRx9px5gIT5BRRuxofs6RGxsLSi6I+Lo1mzYIA3LlPiLa6Qni3Vw2OT6
mg7ydt/+++dBAGrznwIQwUCWdmDWjDNMFxS7M8P0ZdfFZIEVfvx64sHpoWabAkMqzyFeCaehv5Zp
vQYvdK15SV/7/NN0pRK9+566gbPTvBcT6fJu3MxOveLV8zAT4AHnQ58A1BOR1dMM71O9ggTYr1Qu
LN2o8GOHILEu90o/d3qVEthORTNb7mwdEDvuGg8M6BSHBMUiB+zrfpS/BRZdH3pjMRwpD7p4XT9M
6htuYE3qfsj8sTg3v1HJ8sJ90pdh7t6cmCN5H1kMx3vrZRzQJL+CaUtMovCXbrUVNEpztMMInvhy
RADKKKx5ciV253wIiGUHYzoXGavmANqTl6pGWJwr/GhrdpJIZ0jGjQQVuKeKtUUAvyFshMwgZVOy
urnh45x0Aupr5HrT2P6WlXDCs6+gmWGttBLkOzXrmSqWrbDawy/o43T64IHCDDEy7F84ReHjMuOj
DPO5sVJs+7cySD77CwBJYB35G8LNMT3PrqySobu/BqLAaRqqkOz90veBZ+fAOrg3CQA+RezQ8jfL
SHuARLvaAew2zikWk0rZP0HAXNECtEol5lYyTVPLwfnVPONfU8IEbcf8n2K7W7Jvvi9RZb9CFR8D
DYHLcaamdHumOAeJv9F2iK3H72zVxGG9rvIUokp9y6g069MNQ2Vrwo/JyoddRr037oRBHdDCN7eT
tdWul8DCCILC1Lu6eNVlA/6AWyjHlMlFGbSZ79LuyNZte63RTqhSMFzLxQBaRDy4dK5GdPgrw0TK
PX4oqTYcAKR776ZA+BHnDCXpCcQJuR4OY1ixMgwtxTidOm1Z/+zACOgsWLiOp6KTlj+KLIlYmuTw
5TtkyiY2yYTDCRny0KwH8pj3oJ910qL+GYpbJBgdPLD9S3in37Y3d8Il/4kR+imRfttMCkC+VkNr
jAu/7hlU38sbH+/ThNWlC0Qe80aP598fbyqFX5ahKEOzDXAzI7u0yL/I43W8ZQHrgbuEU+j5ctVk
/CVn8kg7x7kBahpBSE141ZF8NqTCZBn2noa0IQotnoE6pfe93JJ03VsJFWijtLjH2SLLn+/MaeH9
eUxAbuplpLCZuYfgbB6Xwah0a7kbGr8KH52EzgJa7eHQsVOdbpacw0ha5KXrqCKpTzuLcr5IR0DH
bU7ZvmPrtyfFcv9Ws5O38V6qRzsi11vIo31N4tCSQz5SY3vcK0yhWfKVGTclfCfEUJWrQiuB0zev
XFfnGAcnpXNP6Ru6q4g8Y0071dSkNycl599dKCgSN4uKGP6yE5sBfr0qH4w10j3sOC0KM5/gkX0B
sYjtd6wmJNkb3KzhAZZ/HFYvpnoU8MZzm5du/udbZd9pJFzyiz0HTHjrluYSfXJ7Pb7V6L9JCMjO
/p00pas/rTiOa4IBCrzHs4jvsy3JtWGUYkbb4QxMGTZgpZqMOZ45nGIdwZ3DbmNup9mFZ6ZOQOjh
FWwn2+ws6iJU7saX7BsVxMe3HjhBx9FFj5IXcmMuenhh/e/cNjvPZewZSHsjTqbtyFS6tanRkU9W
vnsv4da5RJiUHPaD+qeMD5Iyp/xxp0LKy/h3/Z4lQRu8fgYmx3cio5nyctKlBnzIaWVu2xexVDCY
BY9/uiKxvG0jIOvmmy4wN8rYZJaocl0j6ltuupro0vSuyjqoXn1aSMSg/GfXRqtc98ocjA21BCD3
zQATMR5e9N0/HDkI48+oSytiqC8CfV8Ms+1W4RxxKDMdQkinF524Mb4RFrNVMkaXnpJ7GVe3TblA
jrIoVF/pZZrSL+xksUOLxC/VC8mZ9KLZNs4hngD1Eye3UZuAebdGQwj9eEDAepPe6lXEflu0H5Hs
7ktnmU9gPLhbp8wa2THBErEAGviQwL1QWDQgSJn9gy5p5YvsHPBUua9GzCQezCDb57vg/JwLerSo
gFTSGev0TSGHb+XbFKpAwRw1y5B6T3HxxwnMnaKWWWsrQqSla80almY6dfWCzvR6bb64yKWjRhXd
I3l1r9giZorYZgM3x8AwBP1GCRSn7q6B1yHfjylPQAaDVkP8bkXVagM7sOhiaBAUEWrCqvikcHEh
D5fKXyGMGOgr7Bpo9GkC4i8Bb0oNhltrhYwvreVhu5dR3DLb7z3iwhB9GGpUV5QsNjV3NjyXS6hu
u4pmWW82OtAzrsc9TouRhhpxKjwEixA33NPW49tnuHP4oxCo1IhxPvtqxY92DxZD/6ryIqj1CHMn
W+OD3vZE+eWuuzDctMqekz42CcQAIXEIQymNiuHiOk5XQICh6S8NazI7URAvgaPc07UyHkZ2huz0
7bJQOHlVC8gtBW7AfnwZ6/fInjm5+Fdxq0i/b1BRXDPtQl1BkMkMo1N7t9vh5DAvU/QLlNHSk03V
kJjidNqWpkQqTfYc1WVQDbOqbpwcSDl8wPdSf8fUMef65ATAqingWBcVhGcqa76+mYnf9UdCdNua
NPmAtTvdLlZB3TK2UTlQ2KjRK4/vX4yA3bBNnnB7PJnPu30MAxZbBO6Iem4PRkCNZUf2S8lTpTob
TO/UWODTTNRgkxy0k3rf7G8Iw1GCnozVIeB97FytfcQoycKga7ttswZWnqsCDJBAq3lQZIw9APXI
+i98jodwZZmIoQhguXkmgoVR/CFgFPMPwxezvliKUEc08VTCCO7Y6CVsT7SvuddRQfGv2g8kU1Ly
idUHYzOHZ4MrEpS8k9oSZyVwrUw6OwVmPOJy+aUjuJgFWoXn2JV9FNEYwQnYr2zwC+lOL8NBoaJI
vCezfqPcZ+V0ZSBKCaYPRZ5OQkoIy8Uf8AwXhz2SBhUo2WlbhXKCLg4dGSaRiROMlkejtPxjbaaz
NrwBtKbh399RtArQM56N9TQmouYCG9D1ZZoZKfL6m55bILoejAPNfwfMRwPa+4A+G4twNv+Y46TW
y3oSdAPn5o+8DG7D1vKq01t33+TAA1PFn9kfb6PuWe36h2tbqZQ+WVYGHRxqOPxvNaR7d/v3uv55
jLyhE/S74QjjxC4cNjU1ktnK4uvHVXzZBoht1XLAwG+6bRJFWEUvQpcEPFVNY6L/VE6X9wOrDKSP
jy0am/Zk1hiEPrFIGvzR5twTOxO1Ky5n63/4WRwTUtZmn/kpCbY+p9rugd1QtvLmE3z2TP23rNOd
e4ndl3eUf0R2+JwXImpTe8Z9xWkBNE4/KMpJHS3mnef1rz9EZ6GZJqYAERZzO1lh1viyJxxa5VL0
VuCqNTsEPnF977WIMDDFiBVe2yPaQFkHnKFBg4i9R9MMrH7jZ2D1GjlPFsWaJcIGB8pmYfP0vLvM
JBC2cOUkFZtv+MqNh/p94qgbyeKJDk/8qJiKiDIWuVs2SfiqQvksmUCIpZWF1VJRkrwqdSZUkvQ5
xgLqBHxUJyY2Nb8CkU+uJaza236yhCz73wKMIU4oPnMg3DZ0Wo1ish4x2YirQDBq3WrXJ6RBqwWF
HqT562bc/U10ffSAV24kTKjd+vFw3n/qYsn1uL9KA4iv043Bs83CsNvKL8JYDi6Z0K+xrJbVj0xZ
E11VuqzOmxW8QN/ezh4iz2qqNsAQ1axp+nJdkF5oRidVlGT9dbcK3hlL30KoFBg9e2uOZLVYjTHx
L79ChD6XEnElj5yOg7K+UIqhPKQEj+80bkO5CYxLXQ0Uq0Cvz9zef+1K+OKjsenhcFGQHVl9iAHu
o3YpbFg3BYvpOich4EkuRehmcIZNKu98OeOx5q6u6uZ7aA8hjEL1r1yZGTTOUYUP83n8kjOwZBE1
xrivqEv8e/TyK5JNdH3/qrINnE2sw9hfZaW9aWGOFOUQos5MYMIHeWmSwO1P40bIXPRxNdBg2Bmy
3V7NOz9DKSzMOxK/1RGOH3CJ2YYx/w0tIqOi6cH9LS3aV8Xt/XHgZRa+qEky7QdGCEboL4XCwFO9
yNvtWy29MbYsdCAXcSaBnSDuZgAhN9/tXJxHkFj8Ppvrb+EQVPwsYRs6X0PHXzkTNEfmCI0yZUm9
xjnzJ1Z9CylwIGqxO2k/tgoLi8i9itCG3QUHiqBEFXZwND0uECa1tcRMbUHjKtPBaWABX3frzIJl
pjdH9h/LbDIQNwSuoNlp2tuUB8AzVTkrK37Feh3I3cQdTDFveEHYq1IiY7AUMqe+Ur95r16OLBy/
YvqwMEMmqfJhOJ8a22IiYuya5zB140fcs1JY+6qOnINiuwOUqrJzNRw+S1BjrRPGrNz80emQhb8z
yYeVw8DvWcAU7+j4tnp8BGUCJnPsjAclbPsVqkB0WvIuXBcOm4l8I+0d5ICR6CvFWkLj9tKVo0QU
Wt3eGVZsIIWgNsW6kWRxs0IT9xURCQfUfTuaLaBDHoksB/F2AKdR7k20e0Ii6MQrLRG2MvpTaSyb
Kx/DpHOkpOz4Dxn3TKIipa9I2nkUxTJgkrZBp+wLcbF+wUTrjFLG5uP8LKfjy34/9lni0qjA6hQx
Q+SuVOvoLBa4SfMUagfMrOS+oA/CnZgFeDE7Ya5A8y3nNzf0WynqEqcPndQC9h4sRmIyd3ZmkBbU
o7XxEdi//3tMn8c9myc+Td9m1ddenqmzH3THvK7MbgZ5kSUS4dl2WUIxDwTo5YKPLTgOodCM7PRA
HQcCX81IMNErLhLT8M0FcdSeDikVaPgZpFalXSuQNzXhC9nP7Ac6x6rxNPMNnlyUoQ4zsn0WF9DP
Uhh+IUjY0zXwWhFdI2Nzdn06P14o1MXuJ/yVsN283/nX+57TOg9sNFeQSTMLj25uc0RBvnsr1KyC
i3qCs+R9Gvx0A7gqcSslqaaNuKbpuhFFpJQwcg7Ai8LTBGzzNDYSQ/8a9DhLs8q4NilDm54vc0/h
/9oE7pkvgIbupzaaO77nb1mKUJwq7Sh338RhjblXC5A19uxJYIJcpPhfQj2w4I9vdXxvpbSEmPl6
rV27AT2lSThkvS29JMgkdS3nGJJwUelsANTctUJZwYke5AtohLb1CEWwSnHxhCd7DsYfTXfuYSTo
jIBouJSpYyfb2JNfcP1oaQIv4Ao+fmfEKBnEI5daYU+upKYpplAQb6CvgWBdoClZMcxF7hW53bcc
4mPU7fWZfOesKfOOYNUfxh11RvpdC+QUegnpACV2Qq2zDaRGsAZwu5uw5of3l4UB/m3HWqjnHrr4
lPHydyYEaN1gXH+aztLcDcCoxkk44f5oA+jxLVSKd92SvQVtRUIcTbEJYvQRUbI1vGj+E2WeZjfS
ekeMz6+3GSaXlieqvz4gV/lw53cLiCSjIvP63SBo86j7tMhdZnlU9vh/oNb/B/YRCT72Zgfcq3iN
VSJ8KgrUd7hPH0W5aEpAE3zNZs/h/HDbbgWEJ+iUNQwnw/HMew/AV291Xms6q+TvZDdBY4ohrYQK
ymppdFEAzQDUWGiQu2mnXF9ri13+2PvKMsByott/bLU/cnoMZGtgeVOuCxvTzJRuGl8gqAxMM/su
2VE3CVjMbOf3CScBsh8sR5bq/rF6uV/YCrHRR4RRTifAwfSicngkS/4RsIkDxdpql/1Hs6TtPbkG
6IZAYu095n6kWqZwVl2al/0WKvQf283bLiAIXLht6EFyy+iMJgCxgiQI5uVO4LEZaygL2WLloZez
zx8uCV8DhGy/QwaOwJeLVCnmg4AEo1ltRG7vu8ZLNRonDmhqjhJXVlQYNQScFw3eNbOkgqhPizkH
GaQN5NeInr9VO+0esrrxfuNU6Ay8M01A6QEDX40GRTOFZzUNB0hqiFIfHDw46ntSZ7CSiBVIVQdP
m6yb9+U+Klk0qV+x585nh0nBDqIm+MYsrna2BPLRBqPUmF5K8aiaYehAbn/czSYeyTapM4+aWiEB
WKweTphY36TDYAoIRwngdwZW+oOTVTHThPfZ0fLchgEzXatHQdoBv0S0BU1nI3TM1bLL9uKFLZdr
L4FTc/n+jIb1eeCOgRF4TwQAiNITr4NI8u5JypAY5+pZxLKjj9qd4n82AbuGANBcyCCjl71bcz2d
HeBDtxiC628HgjL45iqd/g1OS+TemV4rqnLp8a0kzWhbpFBFEBnmtQZC3lcdimfyJces8EqTGdWw
oHged+jAGrm6YMdySFTCZEFBchH2nxzwDyBAA+gEEgLSjx+gIuclqHKeGc2r0aAmd8hhfDBFNb4l
y2dm5GS/tPsCNXS87Fym/OdvwsPhZGrMTHvNZN859EfdWyzAcrHMiXeBFxRXIdiAasK/QlNNnA9r
ZZ6a57Br5hhHMNPZ/9ZTs1rCGtsiBs3rKtV1NJI/2qsC1ICUgInL12m3NgkumgWIFe0/Bje7UtmD
X4MMbz5Hqml3Xut4//tmYwugHQUey+7ERDaG/OTOEcbh2IkVCom368Q4tpB6ocF7321WuhEEuBiv
xmskrSx0L7UH1FpQvfiQlOg8teqIc87opKKd8cep83n7cuVWcZALvsjip4oZ66/ekFeAJcfFwXnh
YRn7Y9uIce5TVLvWnuMbRcWRwwMQdaItHM7NzDBYefR63Ze6WNe9c7oB5HXXbagRXJmqBDdeVa/l
8Mt71a4YnX29XTvCvA317+a6fR0VDy+231TylB0eMsS7wAPbMRPuiCYb1uFWtz5KenrokZDlczPI
IkSTR2tjT2914u52y14CUmZETwu8/H53w2Hwv47l2DGQgFGnu6D0oEn2eFXXfzzlU1ydL9hUATQ9
5+mPexMFknbyp9oqlNoR6iIh9LvhTgDx2QsjNlew/93wJzvwrs5dGb/Rzd/zVMfwHY/5Z7Oombex
8q4d/15uZN8J+QM9kTOwlYWiNKsUfoLbj3ZbHmAibEuS2W+UbtXafm2ieBpqMrAsflz9on0GYFfc
gwur0ECCJHNbW6EMymXVFQHD13U3zmtacmcbQxdCL/xmrDNSFGteQxSQdLACjw/ocxnM+hkvJJoq
1Ay2oUsPmRdQ9bZNvT5h8ebTmGt/jrGwH0LePgNlmOVDoloB5GSc8A3IvTNilgGGFHFXYt4dmlwA
7u//zeMjVmMHEfsNHw2cOSXU4OKY1jd7OcDwoksE0hUyOHV/7cFUe0Z0+7CryjL+JWTihvs1mzpZ
a1rBPt0m6r1Km8U/H0UW4pfbpUQC/nbhYLON7n5H6maY7XLIre5IUU9sjlD7fmz8HuNIPr3kSeiX
y/uQowxg5zx5x+zpoIhEf6pGgvHLnL1nezwwnqeLDadXZ1r5n7lZXkYngR4IRSJHIjzRBFjQvuHn
0WxV4dsUemVOfr3PXk6R+O7hnIgAKpM5xSHvkVN751TkZKpw1sXwoaqjLRMNt2VgGp697UgbRDy+
jZuzMRWPQYFxZCe6N1pTDjZjwG6M33ZRbV9bv20V0QvCFZiXQIWVXOPQ3vvVKEYSk02mLJ8B5buI
uG04/RLh9liJc6WOPYukhcDaFOGwN4+7XObQM2/iBvq2ReQHK1T0QESeQeBr0nRZFPbFxMFnmUJ8
QIVk32pzPpSx4MfJcXILbiijp56uQH6g+vadBAFC/9I+6q7pVY1F+pGzqqJkV3Iu80IJc+rnZ9tT
Z01o83msT48Kc1iW2x5xPrq7+1X+RmJwA+UySxMtZ25iLNXq3yD+MIaK2DXrgqUbkSKjitebMgit
BAzFgUKHM1tg7c9r+SM9BNHgqC4p60HaY00zJMRxkzXmRlUzFdIUDGWmfVCxd/BkWOLVirj+Kz34
+QFwFQuwxSGJfY+lnjUIsYWQ2Orz62qds80KHv4Y2ea4541Irm+yii6DkK4PLDZAf4aNFGJelhCA
xEkH39zUVvXLeUaQotZbaOWWe6KhkMn5KYe2vMsmdDkL4BSPMu+yJ/lSeom2z8tNo0GeigQmJfDO
MjtbFJDn/vvjRHysJQvaoLfuPGOW+GPgYNb6VJoC8HxESpT/brfuPyjAZInm3lHO6XUYMbJOnt/u
KJLNIodexol+R5JLflOs1njCykSDODj5gnJCSAHQKzpvu6iNNVUkVqOuRKRdf/CfZ6cMixSf4sGq
xdP3jXgAE3NY/vZ+CBsICXqWrKDnwIQ/9RK8BoVPOhXd7aAbVPy659+a1rJmLrn62S8YaRMigCJI
qiRmYLu9Y22dgHV47298Qetnkbgt+l5szzVGDqXa+CEk0RE/GboU37EmB/zUwbVGAJsEFRBOP3Ih
A31Diy7V+hSyJTUOegFg8H4IPFPOiUv1S/Rp2u0QBNbd6RIRKO6Op5jOKET92aeNN6kuF6lTs3Ao
w6oLwrUESyP7sicXJ3smRBI6PSyhNFXvCN12ejNDjpbUWebSpxNfdF//I0vc4yB6j0lhL3jmWdue
ua0hUxNfoD/yHBlpupIJh+SaXBQNFUU4YnyQNMfEtr+89riHoqIsf49WhJ6v4vGPeV3mXoUFPMUA
zOLrQOTdkLz1dGLkarN7Jq1RDhKk7w94c4ENn8TYkaL5Y0H3nijJbwMFsBDQq6cnmhMrdbQloDn8
Sz4C9vNdg6BX0yasasKMBiZILVeQ85RT7wIgzJU51rXLmG3JePT6tndl3zTsaGyEn1oLIRJ6/ayq
tMirXz48soJXGCiZVHpkZeXro+lDLmJWcJR/RBxnL05unigPCZo/5PKL9cI6ePppM/OVy5yvVeqv
E3vfWPHcsSwzvllg3zIqDj7vS7ZHB0BjYfMZK619NXTzBbniNHpCPsUueRV6eZEe/oFA7kERMgZm
gecN0WnDO0BxH6feDQUB+AFzkGUfG/4kbAdfbwPMod90aJMY+PZehfnlwr3+MLQ/5L0HWDrGgQEg
5Slc/4c/V3Lx8UTqtt/gL+L/h34DERyUqp8LC+2k/Gioqz0x0IwBrKd3Zz3FJZ8g/ggwBAnk2Gn3
CrDX7oOFJsCYxWjLKL9GucZIYfyIjfs6QKpBo0FJgcuG7tojw+XX0tba1zFR/lhge9AAD6M/ZX7s
SatV+Cqb9D7fEOST46aMyICE+nOWuG3RJoTYz1BVXOblbuIoHRftk6Q/e7h7WhBBHjKdaOiueMa8
B270bEjVXff8f8wC2TcYyF8vChhg0DKIj1I9s0ywbHrF/coPYvwWhS9qnBeEZIwYw1NqoKUxr/ry
6NJhVawnAQppatVp8OBzyTdnNOHopaFIpU26kWeVV6jtXjzSU1jaBku+fM2YrNvAxHbMIuvM/1RE
O0DmfIBpWODJ9dlrur89MHvZKRgcWqnG8HdPL2iUQXbOey/OegdRBH6/8hpwMytriF1afbNQ5LKe
X8FoO0l1p/lDc5qE0SKZq0MRVGnox9+KPTld1CiZsETDSn6gLRG9aDmoQ2IZn5lCyC3bQeCmNwLg
e+XMeQDSiFWwo3p3hA3n/iN8wSi1kR2e+G+zFWGnoU1XqZbgUlkEFVsHvyRR5KH/MB2WV2DIoYpq
WvA26z3IzXIhTMNaxxzxiySjCfDYVhjevCFlKBxKnEKf5TKYtUqO+V4xg7gBOK9I93/VoPNIapiZ
5QpZIywWQC1Wzydg9JYTNUtSW5f8swqXmEXpgxqItfHBBzIEff8xg6JDaPW7X+iVAIr04K7lZBoA
yH64KVAV+FAgCNcbtSielDlnfch4VjsnsVEuYbHcFqMWK7dcM3yjKd9DUfAnTrm3SFvB+2zpqoZ1
D9aXslDRjsp9rVN2WqP0W9brDtoELFpesqRjmqiSnsB5pIxsoO/JQ/XQDm5CYzcSi+j4zeP2CFGV
xd0AyUsmevybCU6Mi332Q3rxUqeHd0ELmfpj1mTDa/MPC68ykucwf1hy0eobdU5w9HKqIVoxZMw0
WiIOeO4BXT0IZ2gv20ofs3Bu+smZmHNvyF605/Gp4qguUrtRxyKrIIWByEymocgSt7I5UXlvB/wQ
JlP85C099tUMu9KxfvCafGgLD73YTPFpCoiof/OkrESbDQkP0NEuDOGnlvwggZRJqVjokOAWw+BC
6eu78QFPZavWu9Gf+f49E2I8X2FlEzBSKw/2ET3B46EAuM9tr0ePvPzsr+y279aRxO3hFiGN9nML
PQY3sygSD2aZF9wBmFmbI41dlrrac3e6x4eE672E7d+IG8IQOew/e+RwpOA0jvyVYOcgrWxUnIZD
SesbYBYCE0wT0xtiojYgTrPQxTAOYSN3GxoBfrNG7l2S55CaxDngNvGeK6zWRaVEE8DFaVuDTIRP
7GGchfUMLF34F2TTZW96PqD3uja96G2axW8bl8IY+j9boUE1vhtwYwar+D6nQetTxebbe7R11WCW
HCYFwI6ukj4djn36I7oZOgX3BgTJOsT2cpJrBf5VXj7rqDrUCbTCKD5jtBWxER+3gq5gGTCpXFZU
rg5nYasT28YQUBj7hxnCcPXu5aJcE+0lRKGH5viJ6QJezir6qON2B68PHJWn0+EpLSroi9WyXBtn
Kx2EG3B+C3kV31QoSo5R49gaHAnEIumNUhi+joMSANo28fM2+ovrkk79xIIBylvM8xMoAGyAhQwy
XXQukzBLeFI5/ee92Yo5ft42eMC4/QoA2R6jpvFxnzsh5jwkKM36qji3QA+H/jKGSkdGPIgcTESr
/TovB7Xw1yTI73ERBu+njuPWWrJaIQju4B/iXJBBACP/z3sfdEoJamBo4KZ/s93W1K49wgFtfS21
sq3gfUaSLIi+UmN7SXYcCUB0yb+Erg3EIyrQbCz6gAJNeWfqc7mGwS3W1TCW0AMCxCKu26i1oocg
azBpIVelzd5CIpa5f3BvvFECt96g0BDwNNsnEbpEkMYZVmNJjKjxSEvSWZice7exOnc2Sjel4RKg
GRBPCoyJ4k/6tofKIG0m7x1YF7dAyKsWC/JPC0273IVtXdOUqwCoN/nuM6l/tTBRIV9+NAz5Rang
FwiRnvSJvWk1G5AhHuR/Bik+ht9LHrQVjRjhstz0DIwYUQJA69qUYuze+oRyK7JelrK9DvJ8FnWd
TV9qtQOL/ze7R0OhGkpJlv3u6A95K2+SWmTpfQWh+VK4feKOeQnhnQPFpYMiNbu9XTxIeyP2VlEJ
TJ83+FYEHmTqII0zyLDnE+DiN5keA40OQmcwH1BFnzS88YklG3r47uKm04JchBkAfnbg0bWG3W4Q
z7wH3MnvL78BKdfUTqc3KrrEko+VylThU00VTh1OfAQ13cY18IMnu/celQA2akMeFGiynu5EUyDb
NdlZ/VNxkCrurqjLpzzj6hYjtKdkWACB1GIHpmCfRITCSIWEeQ3furuvo4nu6rqDWZ5ip2ikv3cy
bnl9oOlrS9UvP5uQnci+64rIjAiiEvUrQUv6rFSiGeBiRaKIkB1/wPMbkHROzYrDmqAUCj2eZvmg
ZNQkb0YDECMSe31UxFdCqAMUxpOPXILaaoLp8/AcZIeFAc2yercXWgGXv+FBeE62vx7NkrIMRlM7
9fBPhMAKkwsVNszkdMoK4iL63+o5X/pP6bw0MEqQYKOUF59AqmrVeBTUWG1R9Z63u9tWHYFi48Si
1jEGNOCK45Fs6FZCzKiqyOjJ7krfBSXO1ji68YsFH5lFy0m+uhh7cs5HPVQkVUxlbMCvVJireFlh
ldCqsSm5/L/WIfyIauY86E+QQEzMw4DnXQchgfjJ8OltZZjVDji+elLLEcpkFO4pEC1/kOyu3QXD
4QZYZrm2J1H++vcIOD0y/xGxzdA5X+3LUxSd2RBErkLM409Q7MeTKP9g7Nc53vwM19m3YWcO18CW
+gFYsg5huO8NPWRD0m6kQ8Z6qgk9oFzQRh/lPErFlYpjbEVPxdq7pgpRqdACELWP+sk5r0LfrWDv
7ZtAXIEwhfKDHi91VNLcrET4Xqo03blEmga+e9+43EXG0cb0AY83yOjrQ4SWVYUQmNmGknHRGkx0
l4nXh7PZhzY5z9pfeZ38j+AvW23S0XnL1OvNRWSxHZZ28pSz8fXBw1abkbb+n/u6KTSSII0dS7Q5
2LwvK9vEA56SD20lfKFXp61X1E2dJknASjoE5+pe05qq0LLq6uQ6D/B3pHNk9MsI4rMHn/mGpXnH
6qd90e5rt2GDJsMqh1MIO0s35G6o/kJKTf7bXLNDMm8WwQWdgmJOUg8nMlhGYELvLq3D4POirfvJ
1oVEuXDClFYdRLQlPDNdkHLHrucUg+KBdZ57+4yByCTPBFyaSLYewBehTE3H5ci1HdafZWTiyVsx
+4JtJFOyfJde/mCLO84Nsyee8x9Q4A0fP20CG9ImfmT9qWG0ueUOf65TqznINtsvwJHygkPJ8hGC
8fKvrysslAcvYFB+PhtTh2xMnHXcNpRol4R91aqmRIi2jnZSoNzRacm+3VdAqRBscIiI9abRsfuM
hvac+WMAQcwPEfPTknikW8vgcuK249+ZwY3Yku+yvRxVFhJ9j6fr6NsC75SyavX6lSdjI+2aJSvE
GmK6IL4/zE2I8QkPVhIIHJGGqdNF7WUXpTZACwTX2k8LtKJIPToREFdmmgm/qsLSkpA7dVuWBNVO
n4FQUyc/Md0NQtSdJY2VrRPl9VGirfqhKskasnD0FGtw770wr1nhRBjhm2m6HkTZKvAcMCP1BZk+
revuNRAkHKAElMY8ZhSc7dRGvN3FdOcd737N+KrepIhlPJ+M0p1p648iY3KUge5mxBKkxwoW47/w
Q7eSlOP7uJ+CZRwjNri6aTnhwkoYe+ozVP/L0tOL6FSnrCGB3B3DYx01y91W3zAcT0a1P5V2lmcs
8yn6m9BsjdewVDmUfvJP9GDjd6jnY7WkiUmt8uEkcHBL9nTvB/Vygd90zq/uwgJbg2ZmE0g1mHJT
saBAH27jsk2SI5d/f2+3+tU2ULpt8krYM5CaW3IO4FkK045x/RFrB6xWnaB+xkX3mbnuNNnMrQXV
LTnWOjzh0dhGwhBVLp3kOXtEtoKPWorJCz3ae8N+YjlbV5aZPCa2gHgjjrddq74rUtDK4We3A+Y0
NyAPFXHh6yFbi1ZcbeuIlJ1dxAagPgDa+oOhlBwvfPNG/D1mjcStaTtJgaWLv51M4l2uKa9Pkwh7
apDZFQylb5DzTJqOv9fwULptAR2Fmzc7WFpDPbazZMriuwnIxiWmOU0IIysr34V4sqGlNVXSPaEe
n8ocOq7clRZBvvDjEYJtRCdbEpHcDSiGcOin7VmmQjVVGV9PtBwZ16FFe3igAgPHhBQbxV1nbHH7
rIf6HLbIhaGeQfcFTn6KdUxZ00VknU+dfZQN/SaywhuRYTL4cq7KSwRf1oOi1NP2TD57VaWg60ts
4gBRoIVNaEX8kTjL6AtB3b94eEn3XGyvfkZTArLPeSMYAmBW1SOlFbqvG1XKkLHsHmoS1yvmjIdm
KvUphVrRgRMDAvEsrAkZPKpYDr87fSPGKGaNLrNAxqxiu6KPiOnyAXFxGsmOAn4KvppqYqcp7YQ6
1y4ZTBVFk+eFauOiD77rBrzu6Us/JKRCwl9TaZlrlJPQn2j3Hljtiw7EyhO7Zndy1m4h474rRih2
CrdwXL+ZbLCe7+wZVmvR+qm9cwoAnr56+9j1EY2Hqhhnf+h/GZtAUbDVo9vkP8PG0GKYFbFt6z7v
sRWE3bP4ao9vkANly0EN/iOLAS+Ob//VBsWwkVniAy5NddAJGe70TWGaXrtT6Y+A4Gl4UoDlVNCr
j0SZELkzeN4b92+w3Du1MT6PDRUa6EU3AF1tODoM1H2i+RMI6d6sqlLhWwowaSOi4Q0ltbHS7KuE
MXVuhDv65+36FFJVCsHy+PI4b7y5u51d1Lg/+ozukHxY8feBv7enLzhbNDJUPBTr8EVVv4V3nII8
u1nYjXSV99qLgLh7K8cC/CIvxQ4gSeBezG1rzUhKiKIkWDiPUv16k3sCniBsiQil5SolFMdl9V/Y
0g/dXPXw2xRRgtmKADYeesqWvZZ8Wr3QrKXC5Jyx+8x61XV7/Omcksltb0n/+H1Um6s9h/xOOyd+
juc0EagBEhM3xmHOyqt1JSUxtK/d/Vn3dwu31k7hn3PXLVw11duVODG8f+LbVNHy1nB4obPEpDH+
tKDD+8ibnljzuJr+BbrjFskGWpMCno2ypDmzusaxjfwtfLNWLoqyn8SEIFAGc/n2MtXPffsn//Es
qCKzl7zMB/rtRmu5JxC+olmBYKzhnhqDN5jxjPa2eNzeo3ekgl/KlsfhQNJK1Euv4R/VVuh9MgFT
jBVKpDQGki2AwEn0kgykDbxnfOGzFzef57PEYVAAo/vR8SZFpLCEMVUiFMCE/R/Wq+p28V0LRTQK
iV+XW6e+z7OfSmh//wg3NpK6IvX9NLvQ7QstJL41PtEB0k2WNvUNckabGF7+62wl8ilGjE1StLRS
I8ihL3P3A/WDZ1E9qJfifDqafKvB2lG32WkByNBtcSwqAQfAhwitL1WBaLlfBlt1BCZZrWAcLvhG
P+KLs545rZ5E6p27K0Vw++8S5BQRhjvxH7I6SfxL2czR62NRFuMKKktUCZ8Bpj7VnnxkKrHNHdKo
wqChMf06Xd+zx+lmqqzq+yR4Y8JSVtXnv/PCj3dWdgQfcmJGVPXzSjsJP4kUAfuFpFBQQ1hl8cme
5Bb281ZJtlX7ykZ9lRCC3LAxkUp4pVP/oYoftXGAkLJkMbrTrPY4bLyh3gOLZL77m4J/0yJS68sh
UOBuF0ud/yJfwy9waWTkkMZ0BOkhW4yZrtMiN/EJINMjTJfB1TmoQHEW5/vzDpXgsu278dMV5+fu
3ZgZ9WYppDWg0hdrAZ0ZGQXbt+wlxmykWgt2RjUoaS2p51VAnMIpuqBZeT3udMj6OxUUlVinK0I7
YZ916p0/A09czN92AXhGprxmuJOLUjseQHVd2nXX6B3EC1Byen3z+loaEfDGzGR2rJh+S+p5upIz
ZiBtpBikXnBHq4wT4FdD8V8qt7eNEwvJvZrk2efevDEtuRceu4Jh4iH563zzxqKg4rR00lDFYFii
f+H/q0aF7/+i65Gu1WT54YB93QtXaG4vg+bGUZAqlqVgZ5J26Jh5eGcUhZCFl5TLV88qdY9Y1b2j
JzG2mM2ckPMe7pvfG3vz/W2mw1s78rJvTj2cHzEHppa53UJodziNZ6UrYZxpzYaTVETnoxclCBY2
5qbECDqNxPnbpVLfHb1t1AeKxqHKDiyTDdaAYkKLSmLzRVlZvuxliBlwwlGQGjVwMfF1MKKoTdek
S/IXqF8dFZCWQyaLGLuaav1bFefokS40CXBP+mHDum7VKwgA6Z/VagQEnT3uVH77X7TzDweiDH/N
7iYscBA8cN0RXjf27OAHnDLUNz9S/1SqOuiVvYc+vfEam8yVI93Sy2imc1l3+eno7VhjQBoIWMzi
xQFAXV8cw0K7JRNx43R0nd2DZUnXxnvZSnc+diXJGERo6tN7SI7D6tH9eiW5tS85fWQ66dJ0Fvn4
Y7mS51Be2Whbw5JSpHY86J7DIyYaDErzS3Cd8AIHXNzZ0HUAiG1FcpMptZOCs07z8DHvcal2mEXC
TDZeqQKmbUef3xgXZDUkVYPaeY++NZQ3+n9WMi7XaJWI88y2f/ObttJRP6UsBG77ZrQbF3Mo89Mr
l0U3eq+bNjiTqgrJ4iRsDQhtbGPWnRDFZCbG/7be5FS1z7eoKwVSH0OyR5QS6MvKpwoFjIDdu7HH
BVVCBcSrlTZYN3+frQTd9bqbScuJuTTQtKqIzOEVhjB5yO5CHFWJ9bxaDw1LTfUolGflv7WT9t8v
GwkjKhMr2QLjsmnWUEaN2m8sjMLzPUHMWN+ExCbgxrhHWiEjUOAMpMa92VYmiewp1pr88t2BsKXf
03m/bWdcLlf4+lZITgyorAlIcQXRmih2fxrsZEckkoIAeM52ZoVZZR0kLZSoE+T2R/UTSd3an5V+
QWpBL9X1ETRga0QJw2s03jqetOuW/HGYzfFlTHIGZ42ySbaPgx2vkUBtPYfTs45r3j1NJaOT0KI1
BIouKIYco/WIfcVH1h4KQXWNdr94CVo4V/bvnxpzqWVXwyc4d6oJfZmOA2FEHos2P/kMKy/9e6r7
mUGT5SQ9NfHyXYd1tDrZT3dDjdasMZDt4BSrAl9LK9l/3pu8hF9wpalxIF51pvCGV5RoLTM0rlay
hAzt8740ZkClFb8yr5qZHWJFi+zvb2LLiYaQ8qb97sK01+L0pBSe4zafY6+FhkG0RKfS1of1QjAt
oD/5Z5zLpeRd4hSw3j3x8wQGJoGYgie2HPk9sA3VJw2dnO5qt2WCYw43i8dqvxkMPSqmGSssAyaQ
f4plcZ1m/PM1J+TyzRzhs6y/SCozL9FmS+vXEgUAa0QLXDeSM8qVW7fE+MLqhJYSu/++cvC4MCV3
o1e9HnqhHcr82th2PLy6Fv8uiUPpEOY0PGKQk5TMwsJ+ivto8hfl2rAxAZz9uVSZv28lb2gk+QSK
yRilyK/uF+lJLdUDSAnonCIry95igi4gRd/Dub1cQzVd/1PFd8/8K8pQt34naTsJiTmKElAW/ueg
i3r2wgcXGksT3PKeN9YYFNfZV5lIkbluxxOl1/4YcenxTMZidrSS63oApO3sthrnKH5Tnso51wcg
arVCwbu4O/wY5VzynkiOnqb+1+562aDof7ooaDhXrlHbn5t/cgRU+qxXelRFv23sXPQc/osD0eu4
+5NvpbM71lsjZramGFoOTSNDowrBKkMivT2moJqeKQHLF7l0Sd0u+CiCegeL1vYEVTKdgeYcIIc3
jRVfcILoB/2oLHbCzHrzC9EAj3lme6jMokJ6wVEHvIkET7FSZ21oCtyVLnaIpJW+XByIyLxmNyJr
E0Hl9r8HoFaZw2umnVkVs1peRoGMSkBaTgXAnLoWcKnaOr2xzSU8tXYVHdvQFIX61eCH4KPLHPv8
AYd5isRHmXcVqMdJM/yzJJZ4Ck4ZL6Cdkvc6nxtPHYloiyo2/K/DStzEWFJ8CZAxTJqkIYr7sUJ/
UFPeYULEbS9UramBQjRl9sWOT3HlrSviaxrV4P5z8DeppEymSdNjIVswi5uxd9U/gsjo8UWzboM9
82N5Xzg1TeKoVH1wSIZBRn/Bmu5qVnW6cBNjWbm1qqZsOAs3OGd0TtIz9OtoMc0+Y2ZbO3SWtE1G
m5O2Qtc8psXbf14uodqcIiBAGNUgQQyXhbFsOd8U5rCNn+/sG0U8XGJINt614czyo8VAcX+JPG4q
sAB9KUHlpta+9jTPByTlVlDuNZ9O+SfIv77kDmsbSjbEnvTQ9MyROm7bCpQUxLZAxkMR8tE77ZTn
mFHllHqUDnuuHusS8zOSw6rI0xCLWA39VogUzCpBJMFzKXkufli5WMBi9byn5SN7NLQqU2vpiLEN
Mrl1hquayiiMTuyx7slHn1AKjvLkRMmkLDC0vwgAmAeTpD7T6T7TaJxU0U5e+IlTv1wWpLZrW1C0
zqZDBFmmMsiArR+5y9ksHlewv2Mcuqj6arOah50CyOHXLasKvEFFXk8wSfWT8aDQyF+ylunMxAUC
QKiEuSpWirSqqxPve3dKibk1mOCGQC65pFZAWtO+ce+dc6BSvwaDUhpuAXy4hkIrvV7Nqa+RUEdS
rohAPoTUr5p/pOzw+tphH+Sw57chR6WBMxJ1Iq8FBG9qGqhGE6hHO6A+tWS2N77nOGNj/uRFxCFX
4dibGxYiJE4bh7f0Tvhv7UK2fj8TNPpjacgDQbWfxBftKLq0HB7JIsE4biMNdio4Rlp58o97OMgn
s6QOXQccOGl6eUP4tMvVF3Ayum0crm32jnrVLDAWytAjbYK79JXsE+9/uYREfzRwlfRlDEcR/FTv
Aa7AQe2ntQtHkuDkJl95j0svxDnGS2Vm9h0iFTfpwFaxv5Q8CQ2ETgG0MuUHDFYShFMwHGbjCcJg
/zx97ldcTAvJAmEeKw8NZnYJqtwGBUFZcb+ql7MdxS9sUvKGiLZSnh/rc6shYJCjYUfilC+p9L5G
8iNxB0xazBH+tkXA05QpN+CUrFRSsnT6DPMJHGUqtbQlmQlUD/o6XB+Mg6UTpzSY5mXerqzQYucC
hPK9DWG4iw6q3BgTkiSadqQ6JvNbwDwIVR62Ebc/+p4bBNgIRnO9MY5cOI+3CL7yWpxYHhm8mydV
xnqQWhv4mk65Imhx9Roh3UIHRy5gQXaNQI0Chj/umK650B5QTCCZJwbXFq7kODUmsLfCmy37pUwd
ly1+bmFX6/inCSgrBw5kX5duk7yMXQB7SAZxW8mQuMQeM4hvkW57hNjny7D1XhZoywupK95utd/D
086vRFYLXBS/60J3JdPc4XkkpTCZOGDLzq4AXekTK215uNAth7FrNHsJYHV6x1xGRSrSgemM38OG
DNFBNq4fl4b9q2DHJFgVxfCpPTQfBOWbvgf4hh0EUnVDiyxmOirL7wnKZW9ZXVV3FMzTiprn9KX6
0SigIAy1Zb/+Sr3Sr+ceeNP5xD8mpWXqSDel/IfmAMtl8PF/gAB6KQtJkrqsGMtvqRG7HQuhXIw2
O4dy+2mU/yZp20NqLm5uRlpiE+yya3/K4Hxcx9UyuKZEK1e2FCSAafgJuYWgxMSYpU8FZPUC2BTn
0ZoIFHVO7Iyhtd76noSSI9aQJ4BrW17XSpQV6KAmHWZ9GbrPqpuP0ToHS4Kb8jP7mTf1zD61WxKX
W7FGU0XcLRNV/8o1HFIBcy+6Yt5akNJg3hzPRIILf4yAEd2HgRGm4WJfVISZvvarPpmzmuDsuk6I
mmBYJUblBI+xJnoxMXvlfcIjUrIyITCXK93qI/eXviqLZoNs5K8WOtYB2Cc8jRB9OTgnaOVDT6Zv
H21e3XxwmDqfGX7d6Q4XnZUQJij484iL3y6qS/UL2FskwE1lUvPZ0oROCUYkbTZq9TBOzzNfOn1/
g/D7SFaxFIE374KNu8VdueYQn9hAOAiyGHqU5MM2xiUazPbbGtZpYdB+ytXGyncMkCsLAacKOISq
iJyWtSouFHapcyNeQZbuaOgofxKQuO47wKnBkBgwBSKvxUAdiwmb/H+o0fIM/Ko/KjTqMKg4iDWa
56zPG+q0fJjzCPLxlj26l3B8nXK1dGEW5qc8EGy8DipzZS9T2+c/i4GiExzmXNPVE18iIewz6Cy2
TfnNolnnYnex+CWX4D0WeM3sSCpdoqYxA33Wx1wKHwcoyK0QEf+/xZY9+3qcloqDBRc4NrSjKq11
m2vvbR5/6GtuQbi6V1yhHeBzq2wTYQbj3o98SrhzRKKhva9xFlj/evOhZaa3Vo/DWzWWK7QUyAXq
8WktHG+Gag0LVKvv9EupZCU9E9MAaR3dWDZ6JnPvHviXZmQrOmtIEFC1EFle1G8ULP9JT6zR/IBD
W7EzXR1PkdXU9YAGb5qbVZJ7rOUUBH1GDmd/bJa/heuKU4P0Jm7B9sJKWcvPOyzqj8sXmUaXA6dE
s4f7NN0DOqfP0jX++HQ2Z7Tt9K9Kz0OCZO4HY4hycnZU2aqboayQeBIkFEylQjVNsQNi5i8UuTvU
KqRvTYl/baCJ2FwF2EkxalK6OY46woCev+07/JBSYnJRY3fhOGqYN9KIw56uLKXMP5lqIXaxRJvj
tbNkgytsRHJj+pg7XjGVVL4SeJTjAwdSwQ0/E93xX6C770dKiFeqnQsLt5mhgy0RYSg7wT5yj/4n
Ej6R0N4nP6lQICaSUSdqad2PyL0uGYYOeSlVGF0AUAtAEUm+zAjcVmCMlUExAXUUqmk8+DgZZnnp
tDgA1u7Qs9/ccRWq5VLhKSng4CnjK6xg9DvkaFaNEImvUKR9SnLfWT8cYFfow982z+938kzZGwdH
Brt3VcJaDQEacJBdmlIaBaJxDsDm5IlxV4neryw+82u1ir3qSUnNsc4F6MXzXogljBLgxy7DTvnX
6AIRbJ5F/Jkv+xHaZ/78yDfTU8izCLIPPUQDr0LI2LSG5jkAkNuXvfMavMcJGzrMWl6E/V7o1Yl+
34NMUBUli4xAQNh3KpZUeKOUQs72zaLHbj73gV+DqOSouwm8hK9YM3sBPJPUnrZrERlCFJ+E+MY8
hsj3tRJs9Y4yDsZXsu9JmaTj1ba1swvXpXH+eb54FXuRDYxLnE2oNQQHJhCliEwcbS3jmN2Y70Su
Y3PgIy/IfwwaEFJYs+/fPZKcLxHRkHbUv61bDLMEZ8XHNa67A+Gq3TMTGjn/lgMFR+orgui228CF
sxW94Q3KgJ70DBPEaSlqlJzhIm41OqPDJ/CzVTC4vPaqQa3EI5nuUtXLI4elrvsuiGPxvTirmCzN
TPmbFj+MlI7rdqHLSWuI+m6BBaUwdDQHpvLllFTjNF3/8wa+M3/PZK2jhAcyQu2fNmuBfEedY4q9
oBcodDJQenz+KtT+m5MBQXkZtQyhE16bUSoM0l4ygxAE7HKzt4uz2hNMnRnQTmRFJnGKATgyT2b/
w7Rs7zyom7DY4NK6i4MZrf1raNuXn4RqS85cPh+PUKT601b/XR5skETJdiMKrRGciKZa1C7FKDIK
hcacf3G688vLOTQVVUqa9meGKysvbIsrO9H0f3DGQOeaMuBkdp/Uc/MNA2VQH/Kcqri48IeqOGAa
SDgMPrUvuCg7lrJ8BOyZuDh9hnaaUwdghqUD1SvZxPHNOEh9a9dnPT+ecH9+5qyM/XGGZ0cg2nlD
88eExsLLuzhaTd+4DGAFVGuMsj6ZKWh4qrweWBL6ZVd2I+S9B5u2Fek4TIeEIs2CYSYGQtLyQJR0
N1MWqbwmPI/3lJYdZpDV55oBzKT2/vyglitIdwTLm8eKbJnfFxbifJFIVIS/5RNYvxO8w3UD460X
q25q6GJO42VchkVjfnpsOn251FGanJzPDi1lS/a41ePwESF/NnZqlRDhKBaUs8FdbKHBkCzcrY2m
0Bsp8c6XFAnnp3ydK1f/H9LW4uH1ZN2LgmkmIEO5YR9FH6Hzb90DFme9tDaQNVBKBMzvK/WIxLAm
6i1fDyl6PoVr1Ef20VbDto2VMuKYCuYeINusuAioVk2zAidaQxb9TSElbMP4y8pIqxDLpjQa9eIE
ek+LWRFX+PkLZy5UsOnzTyJeN3fC0KC2NYKabwNT4JMsaZYKwZCL2vbyWJsFBxDC3DKsT7eLd20f
zIs+wYlO9z/tGHC+qw2OPZvmp0PcSrS3PQGcn23o9KJHEUO9F/rrLPcoq1bEznlSCYv5/rKC9EM1
cVSBdP/P/DwgyuV7pqZONTBfdI7Q6JPiseEtkwpwb03keCMXEvvf5q1MJstZhbPQtl6QWDWA9EX5
YXaUoshjzpnNqKZmoB6M9RvaYLeXwPel+p6YIg8gbXKqKnC5+5wraMTrhUSuGkZgJ40rE0mf5v0P
KVy5mNuUych2vR0blDpuhBz+gSI+OUj2+0YSm4IFYa77o7d0I/wlP0ryGQdXT9+2aIOE0xb0e6kd
5qZvN4mvgqGGFZ7CZds5RGPeqgVdx5EoDAydfoG4YTfOE2amn6dyG6HWrHxh+7RDHxAUQtf1zXT/
AstqvALPevyRHXiJBsB5oAsozXRAE6F8dbCwKpzbMaO90gbbdzbfyksoF+mR3iYEKSR2+HNGDP60
OXvIJ5xPCnCqAIsccix7uGxbflv8n9wAjvSuKnxZRXv32rI0FrTjcjzOGDaWoerNNPWTFE002iHa
FX02vKJ21C7sbvVnUiN678mny3Lg85uE4WIbE/KhbeX0Q+lYqvh/0w3jlV9c464Yk2KuKTpwb3Ic
91ntkp69fUMdIrsPwRQz7mPtcgdAWcLBL4rMyN/JkLaZKAxPSPZRQkURaFZ8PzbstgjNqfqOOu8Q
90xfcKhcEKOHsQsw1BBw1tQTAJq5mJfimNgQC4OlxuOg0WXsQK6l/5uxycCSOw/ClUs0eli+1FJ9
UoSDstumdobHn8C3hAz0uPDauCNLnC9BFiYO8NKd9SFEV3uJuIwXuj5oZLLWY6pf8aGca9ZZQ3I/
VwVLFJFnlXO0lsG7KrP1IB4LaZTdHJV40A05B3sg2yAez0nZ84msmYXjRnagwx0zK/qJQ3Izi5/L
ZGbYu3Yc+4MpiBTVKX/NSKd3UcOV+CNvb1LICa2FuvoA0DH4YzRCcKgcLStvjQ8sUgcEurqfgBq1
4W6Ee7FMbtLRPh8kMu4LFbPWGCejM8iZh1gN9eydl6krHDcmCJ/PcEWaFdnl1AMz8+lx5bWeLcBP
uCNDmqKHqQPo1nIbWGXxxse/IZtQQqovP2qpztq/TizRUT6VgujcCnBL9bAF+I73pFLIjFwAy/Gu
K8R1ro6QkX/jmHkEXaeoi2zc+OAxRxF/Zr64TRd/ZKel7tpiratNtsIEW/X/2PeKyF0kUCQQmK0O
4lSKHQ7XeAhozsA52LbjleOykVTKB9D9wyN5BZTJLrq8+479RNtFy9ni6LbLO1ybVTpsWog0WGNT
Nx5Gyx+R1X9VQ/8rN9jWFBPP7ThFny5TwjssRcfbWn3hVZRBbLeSvGQVzOIpwsN507taq+yY6q+x
PIxVYUiMkNScLu+7Bvv/JCqymviKmo1Ym6B01gf7ncWswJS4vwnjw9xqwJm/YPNTLJs+yK5yp0yC
jNxp/hpDNNcwn3eok9WjECuqc4fCcZ6DQdZCSi61RsRWnF+Ymvy06/G4ygsrUt2okbjx1V8HXtJt
mYbMCtU5Uhz1tsWd1bK6oBTBShy2hpeoqVjv2RtAS8peRG043jVxT8F65b75ZG9kQMbmfhwWJifp
A/Iyu/m54Xm+ZW0Mozi6H+bbWbBbURFVVS2W7YGX7j1JgegTZftfTnF740a3ZgGI42kK37D98N6u
fEjpAfVvW6Wt4VasnypxUtF+S5IFS3KCk/yQu4Aa3CCsZG/b4hN5s8KGBx8Orfhc1VfYTKsvodln
2PPaFV9caSCoJjSBIFBIJWp0lU9FrNidgIOtD5ramBKVHjkFXD/Oe/gfEWFbFTQSosBy0+Zzn6rH
HwmzRJu+OWVhjGDtzHrF8JUo0RwpmQMVKpp2qai47mnc86ZD/HClTILs73BoQ+CpOgKfr2uAqwH4
k0hkVL5v6UwTHCBmU+BVCHLzfIZ3vQHh7ctmkoTynUtQ1aMHNrE7j0FdmjfCvjU3FzisyRvxILXT
EGFhuQdjWIemWLJJffXHZNvlcj70Li/yDuGUsvWQN4pKPcT3Fr+NMqv74Xj5EjlFCk+RR519faz2
P6HFB0cN8k6mv96uYAI6u6Fhjdw91Lm3D5c33+a9pnk1/fAVjD3CRXV+6rGa1nVtF8qWVALnhmx4
UsAw6HBZHS0VnIOrEMukUB2Ml5P62vnakEkf+el+J/HDbaI+dfhLYvQquARGFraQIivkEFfMr0xt
sYrAzUfJJA5jz8BQtsxK+nGw6ZMp17fDzftqp9m0P2OPX/7N/MQfX/TzQssrjEzOeTgeGUi6pHjL
unPh+B10oOMtT6T5AbTcnoOIQbEPiqwr6Gc/pAKzi4WbEhu9wauxGksKgY6TjPPjdglocIsQbgIL
wIr/jpyhDp53cCRg8fTh1K2qX4j/pvgEUkyTeR4FBxddwt2wKpmAdFLdP33Z0Rw0LV2xWF4vF0EB
Rr8c0sstv9Zk7fcIua8fXs1Q3GYbNnThh2lSt+l1W68esUhTUsl5xLwbn1ocEFl49szthVpmXBCS
MWseUEWScZcutLosuXngfUE8TtML+k8FV675FngPodSpF0kAX3wuyLOLZe5XL/NNIuLcOVIlmRnf
6T4BorKqOks8q2p6Q6AWx+PJ8TZgJRyDbnomQnRpce4AFNMu1FazfsWqMRHCDWLLChZcffNR9uHj
+c4bM7/u1HLGJvDgWXtf/CFm0YyjDSFbCyHYZXgZLsx6+qqOQ8mPU0Nwbg5A2ZgZau73bwqkO5Gd
uhgWF/ADcFPpHzajTpU0IFBBvnkKLEXniZJBOx2lu3CDOdAo3BPQ75UUjrjwkIgbEtE47i9xgPH/
q8jo/g9f6uYAV/EQTU5NrTDoSY9oPJD1garcaO4VmCZ8XvwkS3pxfqxSS4rc1v5cj22P9GOOsoUu
beW9rVREoSIFjtOaNMbkPhib7l3Mq/VzJgTllkmRAuEudIhKzALcMdE9JtW+PFo5lY8PufZXQo32
A1ahkmANHGeDhbIGQsFw/mMhhDZZbeZth2hOrRgIUAtHkcNa1+CrksFs5dTitn/PdNL7ICJ0eQWq
yV7Vhlcj/dW6gnEkkSSuSd8yobxork5Cuwtau526UX4SyCfhe1mrbCfcBS156KZSXt+itJUROgYe
upE0r2gjYMzi4l34QrMrXlnossIlmBFVc8ANXmKHpA/SfRksnxVxLszdwUthVAOY393CJBoxA8Bx
15ZgY8hxyXDc+gec1PshwpBFMw62h8XGUeX6q7oaHcOTm4+dMNYEghI1u83NvqVcwxw+iuY/qhVK
XxasE9inKKEqoepky6Av7i+hN2QTw4JaghGc0fqCb1iH3xX3Op6szYZqDq+sDamxGH+BYMyUHYKb
WN50D5gsAk7XsoKkNhiJ3RX2sPTVgmcAzy3BLLA2Wr1D3WdHmNbTfHIOhcEitJMGJge9F53vvpmS
sKKSatVlDPJP2j3kfX/dCRjO4NXk2OsdWDKdcN6jsSO7TgeWkDKl9fdn09QXK8jOiImR46UX3qsT
tdZfrsfOH5bUOtV5SL48XRJh0U14aIR7fonI5ikCFU9xwkS4hSo7cjJOK0sh+WedMQHYRWZcH7Kb
4Qb/53mfXBcp9eyPQW0LgQl97NKwv/uprQCwe6BJoyB//QgEqNpiU/IupeuBSBm82y9LzreckNMN
zY2qvnu2uGLpN1R2HinXlccbyzYizwul7Ns2NzSosbkjZnEfU5mPzNuKikrM/NNX+rOun4GK2LKI
Y9d8FWPMMzLQ/auVjDudSbZBsfKrDpMyDkxKzCAZNedwVRupR3p2w0EWH+QGADAVziqmbZ8FDlwd
smjnOuwEsKL+7PBY7xrYkQ8Bl4HTwKU9OacG9mW0GrZWeGrg0fcBJ22EqgSG3VzaEQg7ezXndTn/
nh94vETAaXhoDpwWqxtzJuEMH/7aM3Qd/B5YzGuTiMjiOsnZAaiceCAhwV1+jAEy84or8QfarNHh
Z+OK1sqh/CCJOrWkQ43zjqNPQrof3UrOtldqSH0EEEi5A8jH/t6ssVrzsGI7RawOfy1Sb05wpjCo
0YNAlQKV0TV3jCOwWsqEPrls0xlqbZI6lL3B5CSw6Zp4lV81lvcgcwCTJwt7WODb7AFI+G1CVi42
gIEdwTjRYDY0bY6YZiS/LIM34fwiD7kks2eWWAVCCNBeZS46kQc6DEG3nqZA8H5feIFR1uJdKbZ3
5KE4AcJdWEjTZXCZK4qvlgGPNgCbMh5bzGwAf7gWVUBCELl/TmtUvDbgCZRRGDP0/XBSbXFDDkJB
YBa2dsby2Ieoo9Yo9uLIgiUTlotqaO4TnpYG0wblnBcj+My+mCcou1FehtRqWvBHX88rdrCwWKm8
hfzotN4UU/KLZzl1z2CAN8/I2AEeTcCAO0YQ7QPIHZD4rCZjdOfX6MZY5bVg7C4GQHIrufktBJBl
DegWBGIswQYjnWdgZOVL0r0WWBKl3TpxFEKFvAx35hbJz1z4CDVDI1M4GIGFIhWoUxcWgQ5tNS5W
SZSuCJtMiQpqqEOuMvUFjLmv4hVBL7msCpzGsbg+E/xP9mGmstjIlX4Dy7B+ZRRYp1BWPBSy93Tu
GxKIxcYGWilOXgnaA3ylBxObXCdVEMhGh02ahZC3rnFrsGycCkA5V4+f26XRLpIa5y+tejvGT7Ge
3yOnYeqNgTGHdVUY5FKMwov0bQqTw4PgYYkkaQL5SkeN2uSUNSuNiRfjN1FEnWVHcyfBlCOWYaEV
ZAsIhShONEjurxqNIb/7JgYBDE6hrAXFAonBWLhvCrpajuKYZUG03OIyGJ9y8q1mBNUhgRlIEroL
6lslxBHvw41qwYcdrFQQm78AddmG9XpN717Thq1tD08qzlco7MePGHzp2INeqEauj2Pdlk1sPzG0
BGsaB8bcdIPhhHggrkK0EWoSsS48n4HtI0OkIUwwj6Pny3HPOJbTHb4U35I2obbmHsWGqh3DW3eQ
ERZbQMFKXgr3VkUEzmB6Re13rZEuURclqHKrrQo6zSzqRZynSk+HP6olydpkHzLQRUJ11ie9TQXH
XOuAZUs5IMBkV9Z0M5LyWI1krfk0gT1ewk7qhE42L/Z2S19wS/mMOo1QzBoD90I1bYIs+s62aZMO
uzTy3PznuEnhK6YmKlWTgCvyAmzVW8Lv74SjIjyqKPo1H8JuxA81GpEshQyNStj6ZkJasta1EAlI
pDeIc+zyYGuIM7RtYh35kophGFDjAjrC20AJqyjT1y0/qVjGZkFCebDhIkxoI0QgFo77K8Q0bEoD
xgXtXj7U/sJIg4kvqFCTNtECjfuYoQkpjqsj6lGs6obT01lcCcPwinadLHJ6VwKu3ViDsRskJsZD
21eeiDy6cBz8YvEEtePDL/XVQqRIwej3myDc1quaf60sOov+t1omqLcLXRwpNgMH4zUuGAvl6DsU
1Jpo2BkgWCsdK8mXXOzZuCfxXGseaPNBufCn8b1/1b3Xb9fBayXoUO7GPCqi0CkwEkYeuiz26fV1
lZgKQgZAWhglTPTbOI8LvE9AuRxBamBwbBhUgWx/GEl+107INyJMjyVyvpdB+WZiOgDOygKsgydX
ebEV/LsYwRwXAIjvtxzGcqRLGpAULXyMvMihmypwQlTzHWGOAwOmkA5FdVXuL4IXvq9RbWiCcHb6
jsAiH4e5absRDFl8mfFndI/68S8eDefn6RBHeR5XzvEuxkb70Qe2fm71Gac4xdY/pBAh9+iPOLHa
6M4LjocRXOYQaD0l0rRdxfwseGrZ+l8oLiuV/CW8KKya1K7t05IvU7otAd7uJVNyq5eUyr3YtxS+
U9dw8vA2NkQ5wKPnEw4XwCteef4f1ccx1cwEGPOQwziOVE1GY7QHk1bQywGH8HvAekLfrPxOT3Nx
kpuHl6Eu7tUDwG2FJZzSpg/Tx8Md6sbOFnLYyRojyscnnlVtdp8FOfOUs8ZvB0pmfnGVGAar3SAG
Nceoec0Mdrqt4ZrrxZ4Iqj6iYx09oF6JwD1B99rXW14URr0CpLfiQ9/bRtPPyX55P8ARFi64r/EP
5mJ5H4lXluE/ZCLHMdn75vOG0z7wHGKtn4Hyr2rwZmgn9Vz1Gbb6T3QMoKSUSBbLFgwOAN7XmjHR
0Uw4evjZglpNuR1+JhBVQWX/0axkZCkNN5klLNrdAfIoAWUK9vFebXwXfVT2e/uLoTLdQt/SxJeZ
FDmSWL09ghM0V79O4lIlS7KCQD9vDkD0gREncMmZMifQd2ePxqNf/K7HJmHcarP0e0VFKGFgYZS+
C1hHjY8sUZOfRMbvboLH+fDDi/WL2yBX3hqz01GtELbXVVS1z/DDPuPJczJeV7wxtcOOU1a/6MNy
F0jRiF+g65LcNLksk92R9vmr0EbUCTHCl/jHMP/tYkEw3chJITtn6iwCkrQksSpZPMiMbU+uFbzE
luTH3VRTiPpuy8U3IrxSTMtWy6AYUrd1kdZdzAjyN6luxScr9sFiPSU/O+Herp5oMNXz5/taEo5w
YdT7lPQ/THtVUkhkVprTPagRQ6XW2noEuFAiOgHxu71EA1Zpm8EFVRtRIyyT4T6TyxK2INkQlYtp
NEP1duc0/x3V/dXlAmqAzFSCjUwKKNH6HAeRcupAjuE2zUjJzg5QLODdkuDu+bGptzIAUMHiwb8A
QdXi5MyAoE5OTHXKsNFffekUtlOMOUZBrO9oL/+7wSy+aX28NUvWGt/U+OqZHROo/WK8O1sniHss
8y5mi+nwkJ/BCkfZclV55om8UldWEtIBRjvZVrb0L3Zb0uRdBhgEEcpY98YwMJNgeR/Bl/nZ5sMT
uGrMt8VVnrSSmyLz+jG7u8GrYkMZA7fLz58LxqKqXN2sM/eKFzIPQZfoH6hQDD8xUMbIZvOkoVly
syRd1ayq+dchDyos5XoFqkwVCc2WXDSdWofUzCKRiiDu+JXoSnuv1t/YPenPllUGNW1uzf9p7hj5
1He3Zeq7Fjb8i8wEguX+RYyGezAW5WudEQDOnmwV0y2Ij+B/Oq9+RfQP4ctg9zYwg2CB8nXVaSa0
gAP+vMrOl5zXJYLD+c6/1qrqx3dZ9WYN3l83n3mZdJNG8MUUvC2auwFIq4GJzlFZgUZKyyX8L1H+
3yDS4q0NPvPXKbUx4op7/eOM/kX2g/yqO1y6Kvsj0bzpRy60bNH7EjyhsAVIQa2XGjJk5cOs1wnq
Z12ssaljEIqwV3JCGsG6M40NBjqxTTKZozVJx934GmpkrWq7XTwr4bGfxVunZu2msQi0+jMxHRgT
nx3DSKS9KryebRYcFW2mLtrbGXrXquO8ktGdjIW9qrZlAmvYskcJO9mMJG5yRd0c/ysn2rr1giOY
fcpnWA+xYCkxcap0HgLxUUjlLYMls5xEEKuHYUQeYGms8X5l46KUufMT0MQNHiV/LFBQAWHKsxbH
D3rDvnMTXqkOFrQu45WUcT+zXuzjVF3z2wKw3MxxVIueb44QzIZieSuzKoRundiTA55CUiNhB4ve
5VwnMwq2IwDNEB15gSCZrT7XZXbjiO6iCHfA3pcglRQYdu3rbuA2RRGBzGRsLXxOT5Z3SnsVhWuo
78bjGQsP0ea0MzyN+vyYrEuHcP5UbSR+L4EiEMu5DUupmKen/fttJYGJEvf5nUXmDYDtsgwU0gft
Sn8gX8CwwO7roxXAVjfY+AHs/P5MdboV7+9BjL2+FDZ1gemHTponaX/ET2BPYFxe1S/HYUxFVYEL
B4/bpIQDebzlho1778CwO/9bJwm9mt7Dy/0R3uYq09AnTOGClJ3d5lekGBwNqVO+Lraeksi9Y0fK
KOibLdRJffKqQXGMA7AX+DpBnpsJoCfFUcyYWQsbTJ0IM0jHCoMTYlH+4VUAP74TsXkVRCIiSRgk
Ifoy7Mt9YJa6t9Bt6bMp2TLRsVFBvgtd0LOBwBP/73DbPQicWNQMF9OfsfMAvsmwOOeLIQNKgNwy
pArUHR7LWxVbNDo4e2BDITcsE7cK+SSgW/7xi2joII5oPKZDQ3sx7s75vAzSFK5dx+JJo8ino6bF
PGh86Jn3RL3yeDrVX8rSpgoMA2miWosHeJZOqzx9Ff2fe6QTzfx1Ia8Up7YGjC9GReh9zBEQast8
wdgvDG7hLLaK+oyo6KlFbq0gP9xCFnI+zC6sgmBpLuJENFWya9Zs1axqTjL0+k0AJu8+cEezDuif
+nCTZ67z8BdN/SxT4veOFIsxvg8Mt5jxFjw7IOCGA7Y7XQUuVynDR3dZfeONysMDNH/hOfTr39AX
hMQxtqbHbd+L4XBibrV143lOidkFcOa0VnbpM4m+Fbmd8mx9w28gYT20XAq6MlIPZ/o1ryx1o+ao
BXC4yufqSENI/5dZVe+fkAsel6C5f9dMHZyHwMp9lDNzfvw3GYx5uZflWds0HMMkR7uYmvL6WTKv
TzVYxz4x1PAlHJCfAFhnro0PNgEtvAIfkrRb+Cc6AgONLAXgAJmgmoyBKVrhwQPFKZ+p9wx7UnMO
Q2CDtdHW3GQpMN6tvvUExyzczfWP8WPRaGd/f3/5sN6yJUT6H6BEM1Gc7GSltNsLvJqIIKmQt4VT
FC2ig3Y26aIA5JzHJAoWeroEderdalAMgJ04/Tojht0gwwdvipebnTeJy6Y+pnqig7PXBDk5LWGq
x+BHw80OOoc3Yi/mRQbCZDezj0F4mHm+PQLv0NLeGumO8frbi8MwmxqePZM0Du5CFvxC16XZLxkI
+TWesLnJ9m3wfV+pgV7FPbrqZ1wkWM+4MS4ZHs36QZ3/bf7mvtQnEtJeag3/Gtwu0RKZM6JvzO5c
vR/xMdZCLeY7xaY90EemFEy3NeJW/Q1eSFTJDoopaDEKbCozcKqkpQXs31nHOq8aUVn18zmSQFBJ
JexQuFdd4Ppo/Mgd/cGFE9hNWGoywfAfpaCfA3HsV2qRLtXh8RJh9NEDyBbpCltWzRMq8jhzG73w
pnJ65McKR/qH8UbWlq4flMKR/B4w4vRZb67wgj14yuJbs/gvqwPvRBflqsHrSOiTTwcu6WUmQC2k
BzRfYu4QpZ/w+GrvxY0X7mhnxj+zvoPfp9WOPXwBGkQvlRD02pCKJr4PCziGXTZkyqEaBUeTS3xL
t/cgmLSC6EUBaWDIQNsOTo1RTYgFVsH+xgS07eVoX/akUHpr7uZTkJcBroUm+agDBsgSA0XoYR9E
OUSB9kFwo8kOCEZy8F6ZAyj5lil1u4O/xmj91mE3H1XKk2evCJ+Y4W750XJNCiRSE7iaPrJxD3uQ
PWfrj028oop7YY+goSU/QL945xDv/UYy9qDiBOZBo0maaOPTscC7gsRtmF/lh6/1n9lTsu7pmT+5
zUCi+Rtuj93SodCYNQV5vOG4UQ0TzOX0IAtHwg0LD8eEKlHw0HkT6YgrB2Ski7ia+g/aWLeRmtXm
69aCVhX/3b64nz9vEI3FxrIf1SuAfEXNQz7c6ucOI7Ucs7A0FKC5/YtDxNOZw6AWciMjlC7PNCsg
1Ix0krUNspLtj4lPcxUn2qh9UdI0RWooQgDGGiCqD12b7shjsAibRGru+UtDqsSuCE33/b2QihhW
sCIufAjHyE3e8m+3ZAQNHI1ZW31i1O0/iCdPaLv0u4QF0OmUAwj5empfm20Aud9cBhjkz5XNu9/T
VJMuQH6wAph2Eww7o6Rwi0q2JHA1YrkKd2drFU+z61b68eHJ4DH/6P8JAsu4Qw2MERkxhI7yzF1k
GEkKWr7UMDxVbDS/NPq9fg878OBilhAHDfj/osVzKoyaw/eslEFoxH//N1TBX248C4EPZLb22jit
tmF9qP3GRDglkHPUzr2Y1E4P73oCbKkcnZANzj6DqlLMgMz8849FwMvNjtq+0ilAnliU7Ree/GXd
YxJDBeIwE/yiqgAf40T6Sovwiql7LL49UUAg+W6mn3nYGswNVlzPb4F0p82I44Je0cdBKUUNvaWd
MHM6YEVALpXfmPdImyDMAKv4wT/3sIH443xMwqM4zy/axArbbmoYW0blURbWzhrE5mgCP0Xj+7VD
VqGQnyl5x9mR0Ny8n1Sr4WAaX2xvyZ+XwbHn0If1YTVzePhnkaYDDsRL/rE+c+tKguoUVFVRJ7Ut
W494yf5MR/0s3DAs0OGXh/io6L+Snqn/epwagjI+xAdurR9yujzcc58OvVRrznhbTGvtyP0WRzaz
KVhgIIFsx4gud1gW5Xc0COVt71pbUV5oJKFwExuBSOywU41z1BSxFp1b5KY5bEaA7YgxbiEff/WF
tGs1nySzm/ex2RGkWiI7NTPo4+FTB37ckWMrSDsSCvTypppVpjFSeTyi712zfwKg2I7CqoX5EOSN
TXfG3CQ81me4psC9w2y9HwHfocvUlL6Mmgb6kcGuigWpKQeHxQtK3tdiafPld+pgMZs+d/e1SBZr
3V0koHoS/BxlEtdHlHdIn6jOLTvt+dxHwgO1bbfmuiXtQT4oMa16IGRsjhaGwHO0Y0QGfqhDGNMe
tUR9rWqb52+CUloiAV4t7eTjMEdF3nCeUoA4ZSHyZe8H4q+fOg1pOUp8M61d5L3dBKmliG6snRSt
/BIRGMiZsHV9WZZwkskJWJ3cYuC5FDp3cQ+GJefei207FMxhdbAzDAp8oRUUoqUhTVbdy+z6u3Kr
K/j/N2wexXCV+32DyjHEMsiicgWURxIxn4RRN+qqziGPvEzAoAoaM8MU3cveI44zhYtZAopQ1fQx
W0irYyzcmlHQjUN6+PwIiBHVcgNtVEnqi2RVeQuYQCQGvdY+D2eXKcs0yO0OIrteEHaC+bqxJHnj
FssDk28gw78dZm5wDv+h3Bsi5DluGtZxjcxqxxI78AbCuZob7vOqJ7xqevc9MFcW++0qH4FTkTrf
9dpzZFAszOM8xaWv3Mf77PsBueAfsMhPJo1qpZLk8fp2beg0BMbyzTyDe0ErrxP0DCxBeI2+V+2U
RAswlbPyT8psT6xQbpq8ejTGz/ckAYzw8a9JPoPYVN2RU9HMugT4SRPUbSerCylWop77R7PQ1D/8
W2uvBGEEuG6yH2Hixkpjr1sWyvlEWr92Uk6/Ivw+H9RfIMFyXHgeRRxP1EIx/VPU7kHHHJtNGUgt
L1ApgL2j/BkcWE33GhGN63tmbITPvYpq9iQb6Yeq5srHyh1DKSq5g2yGQ7evtXw9C0oNdsWWmtKI
z7QiBPgEgO3Oo2c9s8UCVrlWrlLjt+2fMoZJeAdB964oaBOhN7BtQ1WwFgtAcTXlObDM+pnV4E2w
jNsRKb5W+QHWZEEIAL5TGyhApovthfAduyoj7Aooi3x/AM5bb6pwpi5Bd6qbOfqap+MvG3YfVyMz
ZU+inDY85uRL5H4frpC3lnP60ul7GNJSUJmieypt+3octsq0ZLQ6oQexmuHZjqYsi7TjmNOi68X+
yPfb62LIR6RmF7NL+trh3s7qYOeu4p7umlyExZg14zb7lDTQdV0A14WZeYjCR5ieKC6MIVe1fDu0
+ynYKXTO66XecCdbvgEL/jGpsR6UlNUx4T1F9dbRY5X4HgAlOqKlI14OFf+Mlj3SNeQlxvQwDFbE
+DH+GiPdYPhnIriTve30nMMOPEKkwH9Sgi39hXMeyLkr5xQKid8F070JxqPOZF/ikFt2XPHYQNPC
nT6S2IIu9zxwwvR3/BvBWRYWGCcwpXaMOfTFmTOGDv9mJXgp7Ifeg6JrZkAfAbPqZ9T+96L7h25J
H+Jn7IIeEZYgPFfpnZO/zUT+R+c6fljRsSkUQmYj8dsmcBKZI4twEukFktLZ626VBViHZXSr73K4
iA75D+Qx+yd3QjMQ+LA45etlgzECZ4/z59p/fKkyU7v8LLQ0UGFxl0/McD/n+py8BeFfoPc9DZWV
WdRLpqlbHRrsWlFMsD2Ylv0IsH+D8SjRgYWw6UDUv0Pej7v6dm4Z4zOqNeIa/96vP5lqeXTjX/jg
47A15MKd8xJijNNYC4Xw1XowucaNeryGf1mTCGYXXxvirHh5tGPk5sGjsNii1C4rriAfF0fnYrfh
VMDYUEJ6kr2cTwxWAZqxTe9uj92xrBgZWdQk70z3aFVD73PNyqyj+lMJTzp5mGuPrPt+hRUV54I6
1v+FWvpDBPT2IdxuEKFb+sBmkLC9d3Bh/yrY1pAXTZHPc7Cypukd2T457tXxn4cpSVAGKuV/BG67
Yr+norzbgmYCLGGY/w2ZQMBHfvGhnM4R4nkDUDhRNzSP8v/OVhnHpPXCu+cDj+StkYsry8JSABb8
x8UIo00vMTDEDKbqzM1ZcA4fbAhCa9kAAY3xOwYLsKATa/LPalIMRZ0NzF/Zga0RrtSIK9F+ifjZ
j7U64KQ7i+JELOf91tcxr7qCkt29Jgj/RODx6fEmbfhh5SFpiAuXdBsjIuDcf58rK6CkqCAv6LwD
nvDW16k8ZUg+fm3N7VLbiq9FRwrixsHtUrQhlelJmrRVUwC3UzCzwmyezQTNbh8RDaRTyuM82aeD
aznPAuuSd6Cxv+TfYhm+9LQdARsCoPgDhJVTAsfuZYQowlNUl7/qAr0kvzHDFvUspUNsd5MJvs+x
NWpyBd6wF4yDZQI3rdAu6qMYb+TVRXaPpq4Hlx2dlV5igLcfx4yRuTj738I8F+epx+KWWmqe1Ngy
Qc6hCauoqFI/KDFvh9djRpE9p/n9ltcIHjnML/P+b6aMUbHx0RbU3qru4DD74VqCREm6IAQklpTY
qQdyulHVC4osozQX/JM3CEd6Iz0ZRcv0Jb20Ww0aXy4VDLTW1ETDdFUfvGF//Wxi/XofkKDAp3o5
0ngriQCB/8sdguTf/CahaCErfydMIpRu+25YZAe94hAaTD4ErRfCIzYkTSoGk5WHoqONxZlES4Qk
OxCXeWStaNGbpPBbvO0cY9ZwzQWmdTXZSzjO4r4tRiGQM/hp2uNtDxOBvLaKBNIV8D/sF1wW0or/
MtD68DxLxdIYlAqyJL/zSS2VCKfDJk5VU3PPnbSrZQAzb6qjbnr66kPA8DVj8e6Sq7vh16dWUKEn
hr1Zrihtq9grdDqQdPqaluPMM7knNBLDdo1ntXXj3GED9QuWF8VYJ9x0PxzBv4R+WfxQBhaXMQFr
HK630Y54s8hDR6eUNsCk3WIjSLU7jMYyVhyhVa538wx8/zDipCxki045EnpDg45LYgiIUz6QGqDj
Tc60WumFFJPbwZdG+tuYddhcT0IvEyN9GZjFK60zYv31hMQxFBtwKCY828ldbgmlgH3xez+4YQ4L
ZQOegoVt6u4ISB0a8UtErEKP0Dp3IGplRj7aLDdSM68PjGk9weRrmMzTYQxoJ82lpqth5Tq8dWiD
9sokpbEwdCOS4387WO401s2kXUp1yNKbUb83RJgwam3+2p1DXfeXE/bI4b8yZWZRnfDwRRbXemCN
zUcTwMoYYVv3C3VxQHaNfZ62tRwnQmvMEeCGIjdAoNu+mCt/3H5kt8edfsIrxDlFK2EZnXuH8uKE
aPL5RJYhRAFV8TqDuiQRftj3x+9Gh5wk7+4wsA934dJcfP+2kBGuXvRDHSaFW97AsNZ/J/1yIccn
EJ3gayiV+bdoQ5J+keX3GK4l0xT1l0GtlFbU4ZHBEETYHomq4/KOuFyVcNmp/UZStPqnBMr8YxNG
q3HB7bdqI9IxvOyIhwEqMtimg5F13T8/QaeuK5pe4DakqYin0bf+M/W57qaO4NXvVD40eTpLzER6
gccvTTYTn7+74vjdJSfhVmyB1VimDVXrjlDoErNHXAkzJW2/pbSWmqtOZUu1VAzBv+67Eg/93KvF
hFMyLc4irJOk5Py+55DNX++dKKUrceCVnmWgq/Ss9wQ/b2twxlkjKwVVSxtAEKu/GyQdGjG0fDVO
9l52TtLgbsjVrvnRplHLDoVZ2RTj8g1L1Ck3yTJ5gUN4KP65x86Zz1bVxeiNOFJQVZWVkZT6PM+b
4vAmBz2U43Oi3p5XsBgecn2f6+D58HPkFV2Dvx08ph3CMSDDnd1HJSC0aSIQTgUVIngZ9RnNLD1E
0jVI8GB66+CllEOnk89jqZ2D0ox2dUWchwlhX9lYysey28rvFJnjiMQJcm1ICBY9v5hwJAAct6A+
EfQa/T7uf56hu8I0OreIxVTnqn+5hMhctyAD6aCSk/mYzYOy3n/CWu7tP6lZ03a+LTnyFIhQ9G2I
ojImadj2zE20Y1yvTQBHpBTKfSzSZp5HncBK8cLLINu8zHHRpnO9NTXtAvWzMFWAaREe7QQ+Y24p
0ptJupJwZiXndiX/VXXwBio6ML/rFYs1aNy9E+G3fuKLeC6jnBu8LLdL+oG5GCvucqBbqg71VsYx
i26aE+BWI8bzucg5x5DmY6eRXvc4mURQTN9gQZXwjyc8y+SOtkY4Rp1ppFImBaPDoSwjFlk+BN5J
zgrYg8WpOHTpbAwG/UwPgQJormDSN/X/WXRsN5mkC4N9J60La4UgzhVVe/8Vod/UhmHlevGlgjBr
ZhTNS4xBW+dNYek/3r20HKW/CLm6xlLq26m6EY010AcH/aRW5M0VMYmBkilB26wDxyhjsytl2p20
/fo0JR/JwqBisozc1jeXb2bf0ZrTJKjcd4B8Mw/KrS/UK6YTBpwXVrRT8co8OCCPVs1BMHK68M9r
1ZUbgChUwKy4pJvzk0qDzVxUgCaQLSllzbXzGYGTpDWDPuwlDRcUGFvm0zoBIquGU1ML67a3E6bf
sZ2AoyW5Hc1h+LmE1/qufH9REI0AdcsG5uDZs21Yhk2zAI9/WafFPUkOLhxA7rrqiEWc9FXJruFD
IaVHx7d2Ee4mX6Mrbf3dVfMRoq/0+ftCVzJJTk6qwlGLtVCJgbB3EhAZTqNpCAqbwl9pKfMzkrvq
Ej3xylg7fL3m68wTqsjMEprwFMVh9qcmxEkdC3eAWiINnqUCdQwX+Q16fUTIklH6cMWAq6Og6Xhj
jd09KM/wQcJnR2CSzonGS8sYiN02AsoV6GDfNJud9zsloojBrV0TE6eEbOunpewPRTqzbaMjy/93
FoGHP/uCfBtwBlZWpbRsU+epvztKGmJcrXzc/0ioa0q7eoFoteIfpi/yxbA32zrmy+pmaNJuD/lB
1vXSI0NdTX2xt8RQheNmmy+DToahubts4eDJSvNyK9U7Z6X0RpOFYeTWfVVDfsMPdvGt/B/eGCpX
+tpZFu4hR/Nbz25v6cPbndxVjdOzdOu1H0WlS/+fxgwUDendE8HtDM1efoRj/sscSePOmt+1jv8o
GQY1Il3GwWVc2mX80aJ/L0WKUGS38pRcazyCSlQy406mj9Mb4GNueFg+DZWWz5o7S0DtMB/icLFA
F/wiEWDtQAuLsfdUB/oVkaCyiVG/A3F8Ot0Wd8nBvvC58IiM3qQbzWo9z3HIXibJmzqkoyIFCSe9
0oCj/f/dXaMnf3Vy7448+a9goSIahb8O4u8uh7qouwwqA+A86vJVuPdpeBH4grVK6GBjqPjPVml9
dPPBM751vj7Ww+mUXMDGLhiuNE18OqiguLa2dcqoLds7jef2O7KGPp2/o1k7yUYmeBFBs+2ObkSO
1/vsPv8fZYmxvYHO1Scu7T9S3FWtyEXd3mQkMLP4Odu+sdj0u8QNS+rDmzoZO3RM9OajfJpokZJu
QbJBYeyElmH0wVPIKY99ZRvB/0nCe0KiG2Uagpq2c4TYdaHiGAnLy0SWo8c+xq3KpG478sM5EQYG
GQzcWzSs1QvIPZY3cYlulxKFc6Bm3L8+t1/dRYXZwcoCJbB1iXzsqPtld5NDR0g4W03rPN9yLyGo
/VT8xhYCfA4TMSeZ2kfa+RbyItXCmVUqzktsVBXVcoYtVTNN8gXlDRDsNm3K3/iudQdNF8hVkSTk
+bz5sOemybyqp7aCtwc5Ru4uVITGX2b8F8yzaNi9OC2MCPOWD219UnvJb3F2gS31apAk89sF6BtJ
UZBl4r1+UBoyWrrvTecnWkFaYAm1rgDspgD24BAj9nfrYoJW+o/aXXueohgcClUr3a2hdXvij92h
6xpcVChyqTuXZupmZfRa1GpvlPc+Yjs7z46AN4kyHi1dXzbfCzWb26lGZ5nSNnMB4lNZPqfzsKbM
palvTS4zvRNWCr0V0GChyi21uREfG8tmXVxyCMemHE4lSPVOshMu2zhidGJkMLJOeO4mnkMyrHcM
ONHqhlEnhE3z9IaSi29ca+ghOwM5fTTel1iMoOcg+fIsPi2C3WMM+01Cfr1X+AK0lPkc1tMWKwns
A7I+Gxw77qJ6UxA42q997cUZDC2qFyXbdWADkhB/I4aBjUshGed63wOL7BF3htL1iwsYfqTeaN1v
6fGGDLj0d4M2kYGehP/R2QErwbAHpq6rkAbo2F9r9stCc8oU5CBbihWiKmwvCG4YDQS18Egodayg
T1XF3xzK9gVPedrvp4WRz0qjOaTsNyF1sZG8qZkTWOz/5YF5s4fOOGP7n7iPsw5Zzn/Y/OqUI6jG
avVQPDMus5zlNMEOvSaWJQNBBGnjG665HrEqC2TJjynpupvkP6lKxfpGJ0+u7hg8RBtFQBf8LimD
WhNHKuwyj/8DZK48za0kofW1RgVmQpnA5/9yMxoVl7CUkqegBLg8tqK4MKzgBzBngAe5kTYltkm7
Nz4FVkqaMbepcohHLSq+VRX3KTg6CgAgRBD+4IpqOsprUvBS9Isf6ij6J9PsMxMm7M649dE1RABU
Qdif/KInt9sEueocSE8ioYqr7mC0e3fcWeTxEUbac6gCHsi4NAVhLZBI7WcI8jGvGBpCOCRu4/Ax
jiJtBcCuouJmg/McTtV26nSL5n4RdZobU40U2SMf+sc79P4bvlQBfCYLcPeAK3aoFWKoeHfH4NKH
AEdD2JPMqxQjDrZbhU3BqdotUQ/uPUdH2mbQKlaRU4hwAFks/hSTIPV2gJ3ljYkHLlD2pFBo+xjN
e5MRSvUtnZNzEOCMQ+jBDy5NWtHLo5bnp0YkNavmbsXUW93uQICtxYX2NAY1Lgmow+ruNroIhDLN
t+x3tiNWuBepRaV6BP/uJ3FpqeUCxCL65/MdteGHz3yGOmvVpZo7S4OgVS7sTuAJVqdNYh57YyYF
eqlL4YZ0xLHl+UyXPN8UmHvwajvuhNklEEHynELcyZK/02nCpbcRVv3zjBnmiucBPZWFAb2CDn/u
z3gv3cKx9l+H5qvw3MDO08ACoU7w1j2wR14138HcIejtjDaU8KSrpqvdWSEXMEvtCXMux567wTPI
sSwbvT7OUq4eBmFVLq7VbsZrjpAyna+UzFLBd50gzZRTpI9nf2qjp/ut/7iSM4o4m18mJuZD8e2A
18pjgzwfYK4F6QQ/l/Uy7ly5B0e309nTQfkTzAN3bXT9TCa11Wq0otqPhgqEW24Y8cfv92ihi80W
RNvPF5A6eRi7njuTt3OUBQwOgwdgfoqKHp+ecoDcDWsTXtIzQhWFE4lJ+KyCYXefIkM2VbNc2+Aw
jua/0m0MEpdvzCWaW/DDFKXIN2sT+OMJdFOWqIPTXaiy3D/ZyHxEjT+9S8Jz5BnA4IusfH7DltyJ
v7oxNPBwGxAOYVKgXRJmc8cQiewm7ifh2TUv4P6qvX59tXN6n83XwXm/GdF9181h9lV2GaEtVgx7
7SdyGN/D0a+ZGpE+eHKEKFg+LJWPEAwkbsjotNRPns1E+6O42mAGNLGHLa0cZDtjtq8tDXfkF5Xd
3OLbR9YnZFBR3MTX/+gWu6vt24jTGWp6t95wbUftVhg0DSRRG1diW4ynTVNjplb8tVxiJuxMJA1s
s8++U34251cwU5RrC17+VoLlj71v9MTkuXNZ+R9/smiMUF633k1WqocI0ftwpAVRIMVt888DUXm6
jgDlgOLqiQAJMuzCWZ3cpZIt4Q6Jpdj5bY6pCg4ixI6d4lbp2fnqppY+WqbimEAhzSkddzEM0YDz
JJFxq2A1Kp3owJlMErmWACw6GkQlfLRst2W3FhhyMqzYbHmTXVGEZofC3WWbKMNax4ZQzLETIaIw
h7JK5dDGPeptli2CdLf62oOH5mVeVY0euq4z1I6JlgxaVplOZorZBRCQbAFlUgbS8gnx/TSicgRY
5nWirXTRyga/A46q2ovKgPh/pr3R2l8dM1tYTmkBQhP9DiiUAiLBymp7i3y7ScTkfv5QwD3Vc6Sf
FEKBbnz/JjJI/2VB5u5CXG1evVjTceS0jagJaMjCUNcGLZYOnZzcroRSDQy+2rMm33T0ECHfpLt5
8rVviwmPltCbshBhpGGrYZXAm9kyvAKvUXYUfAMb4IrWyGtQDZhZ98IZMuUq1LcjwmcMd07hmf+G
hIV+Sa0kLllxs8M/62MDtlxFJkTJt5eLiX0hP2PwXJCnEglbUhsd68KUAaF3f6U2UnqqGaVW0D5R
YpZQTv2RA+SwjniOCzIgg/TEEfO7H+ZSj55YNwCuHsXYJiVCDPf1yO4g03ZEk7p2JdAytGsUWIoT
8gK5ao0zpUdHEYILFCZuDMRP5rhUSLjrkiiwAk1Q8RK0TzCd/3/RJBxhwBNo7uLwypW8lmeU0Mqn
dju1GTojVtPaIuAei6dkAhj5HZhGcB/hft8kc3dXmkFKWzEsRAPNnyOfAH3lt+ui0UrSqIj8oXCa
Ne27YMb0GASR0v4Y8DNElQLv+DXjAf+l761du5VL3aBLlxpHhnOdfvPY4KxJ6jgUggTKnTR7g9p4
IZ7H0VJ6OrludAd2ldN3TOdQ1xfNOOlQugff3lG8fEWJe9P8AJE67VIjuaHgZVc0NL59PYIoE2bF
CODV/e83l6y5FIBcwW9187hSy6pfAxSTAdLSM+JkXR8ghXtug98QXcoobO7NxnybguWI5c6EWMGb
cD4As7BXpSEmpagfNKJgZZlycKibZdsHe3tvS62TnxsvVR8IM48gP3ZpodhGXS9LXgxYrIPER1yi
irFKuvV0/JxIaQDAQlhsNyKKQIwGLKldmax42xK37wIHyQ/P9QBIGCbg4eF69XKoBW19SvmJBHpd
YLM/BhjEllrBGxS7fH2JZTFxkhb/wPZpbV2VZxKPU7vda9XkndIlQCILAkJVMdc0/HVZzAaUw3Kn
w8lLRSHqmw5HO7V0Y7+Ud9WIzOTWxu+gDNhJNUor6Di6u9uh18YBeYP1DoI52biSw3Co3T3xR/y4
8FtOXnWHwxAgQmrO82KVK4RxOFhVwS4DM3iv3CGAy1csV86O1YS1T3cP6WrjAA6U8cCDmP1QvWyq
sHrBU5EJg96bGbOr40snmXKy45afVR+MwU8tT+19JeH/iMJc3yEbqaWYZFZs+R4dz2A4sHNdnefa
4RfR1HUJMsC0u/DXHHrNtJqR+DBXw6EYRYv50UYB6jRe0ukAap3HiP8DniITPPGVjkIS1o9BlSvj
saJaBA34EcFdeegELCeW7f08Ya/os+YUrLq9RS7feVcNZLx3UR3Ny2C/3hQA78xxZHU3zUxyreV7
0xFBysEbOu8lBAbrx/WAHrGbbSgOnO5Yb9apgg77AhEqwV8WzWNCmnYGRHccpFeb+g9FNd2kFMVP
rxvlJWJ7g+UbyImdC1x46mfm7Oj+zxPH3m/D7Y0BVQsVu+w8BuRC+3Z7rVwtyl7LIbmqgFF+vJqs
AMP81Kb3HHrQOBQY/PYM/Ii3D/RhlwQOAoCSreDRy4Povp5X630WsnoB+jHTIoFOEe2ZZVu5XLSG
UyNey3LmjdToXrZKSR/8F2Y8fh5hvT806NO0KYmCts6WHme5FV0rGpxojLQKw6pzJe3E6/JgcIcM
b8D6FI99dOin9IuqAvX25N69a/FhirKdomARZ5XjTvKdAEB6aQ++pJ3kR/FpsACWG1m8VaI2GtDL
s4SZ507wuheE7xvL5Yo0Em464rQznzghPaL199NCJbaRt6cbSJcIgNA1OFaqlpkR4mcWOgWfm9dD
F/UV1Roi8gbbQ+Xc/NNEU1FeevvTzroDpQAHV91foti+3miGVQLnMQvlGjaWEk++BJlnTln8Vqu/
Q82ItijIXpqMC0V4SS81fLvYk+bcmRHIuxRW9L7sstlaCYXk4IPybQWCA/wUV8jYAwbTtFuPJxtb
15LWYgpuGBdt0VmL3MBUWDGAb3/nnmvg2HE1qMJwhMD49IncJhPsOpMfEgeZcmesvLW+ds5H0wpY
Ai2UgMfp2y6t3WUdid5j93yE8qGbeVpc0EWHoF8k1QIYITT51S6AmR2kfRHiPvcrzymTb04QBIPw
qTcd+1cdu/K6vnS2oux8MDYj1KCFWQwtx6PVRNcLd5VkM7GccVLz9IHx+eHFepB6s5OyaWfLCli5
JxffhEME/kT6FZIXybAvgYfZiX4c9zTHN6IycCfiCX7UjCx/u6AT7ZvT5rWRg74UwqVKIx6ULupq
5QcIcwP5tuOAyiS4KP72Krc1momqPnlxBRVnFey2PqdUmNjyYKvXN6nzKOPIHEcnoDWYq0uoQarP
Cv1nrRT1PkIHEm97vfRFbL7YdZeQZ5rbOAgUQ3C7iMSdYBBgX9uo0dCJVf1aHZNj4zcYlOouUR1T
4n78luolYDpFMkyUYwtSaREXr6As8f9tHx4duYS9X6AvaW4ZWyLTP5+FWz/JKTS5butNJzyOnW89
Gcw2yEOAemmciz2u4gyqrHz7HkAbxk6Zg80nflGoyEp7BMxbbHgOHcv/qjr5MNCWhIzdyUHjDmql
JxUgmoIlftfxsZqcRYthubEf0G/rTGtnv4cfL5xXZmpvTfhNT+3vg2yTLfjTGsnje0uI77Op8xYc
clPHeYjLT7OdvthXY3SF4PUEHTyutb6RoqqSE35GRAXK5B+OlIdgx37YqEc16TWXWsNZ8omX/BBG
TS0RfvT5GwsfOee9q4zxaA2Kipppv131NjIAhhPQapj+yOI8NcmPW7SxSxDrNDJ0JALJphMUguyV
S58DgDt+sd5FtdTL51HSMN5kB4PyGjXSs2dkdMh65syaON9uu9puQnK1Z6bDYyuJLbl10kwSlk+u
zQpUj3JBAsP7Ol4mqeHINHuP5u0tsVnMSl40EiKOR1q9OtnnhcXqBX5z88Bn+b7lZFfh2p1VlVyA
0lRMqw3evf7oE5CCumOLReYZB9a2eTn3tQOn7tJ1CBEh66aFLvsv7+t+Wv9WKHVrlBZ3txvkPKl3
NhvqKOi5Rxe43bCuT3H1B02kjKqDptpwG8cPEnvHqqaHoXqznDLtyAwXEYqEbJFlR/q+jy+5gq2s
/OYT4zZBWYITZ7MUSYrqREcZ5unN2MHRzYxIFIZKrhAWdpJOh9Zfg3XDnVOOuDU1I66t88sN+idO
SNTxgACYYN8lI0L3brvnZ1z8u4DE5BMINdmUTaCCh7eQkMnKV/hLw2a3e78O9hhKMlNCVeu/aczd
qw2qWvmKmK1F2SmxoMLzTwtEF8FbfDeYQGt1J5pQVssQG76KbnYpZrJg0MzRiI8bmBSdjeu4im2o
MXiwz+Fgk6TTYEcVp6mm6/8JC8d+lD5MozmSJwX/BUzEpvNWkjTDUu8a5jqvsgAfYDoCs4b7FrDs
CR9XLWoe9+5xOQIJVUtvhAiL3WlPiVjQ55UujXjYZlzDSpdYHQ5A9klqXjI/JIQW2dRQaW3UZZ1W
xQadoWLBmi2EENWyRSU63JUoNAiAMpLbrWj2NlRQ5UtbcaBJ3CLpRDbsms8uiaob+t0weeXWxJja
ZPYJgf4KwmwEh/e08k/CjnPXFZvwNsooY2ecVv9KPjKHbK94O1gQg6s7gQMgQ4tWKkaCxb8Sh24n
c0f4WVSTUNQQ7WJ8hykru/N3hTacdSrFg/6S+SdFaOU5WQ33bI0RcOXHo7ta76FLBWEmnvecbihH
ONFhmJ8iujak8Aga6RhAx9OjNJhwW4MHX1TF4ldemA98K+fBUrLF9OyckUycINFbF2ohD6NrNucJ
wJcN5BKB/Ec2PJuQzXBBjqqBV0bSQcTVCW7x0T4eS24A+poqadqHZR8kjdV4metX8vOfV1wlEkNy
SnQuWbNMrNMlUk4Zo6k8PVc5IpygrfPOTygCSmjP60+6iX72t4Ly9IzRTfu0jvVAfLyrl/Niya15
gpe02GT5fKF0CRpCh9U2oHZ683dhkPoFT+iZKjDzZyr1/hl6eiTVMmbGeehq7iKGsROA04QjIDMt
W/I4sGrFziG1o9Zi+usTT0Hh0vMaF8C+CJxZiYdxXfxMAOJYw6G0p0ZD+3L8iOeK6h4rH3Y3c+3R
8h/HdQ9l5uJeOp9Y06JOLNvHwlYLAUXYOvCkzA1Aw1+U7UJNUsfpM6pUCfcKhZbDA0M6BFFUch1g
HyG32CbEQN4rckAqUHm2v4v5CsBHaqvQ2MkPaLFyIIiC0Sr9elhaNyaF3zEWYZrhljOWBPnfumCp
BLldFBSYHEMurfYfXs14+r6sl6772dk2KQgEQei8q2qn8XQX5WnTeUmQ19uNXqM1QU+Nl2BEM5GU
f0z/UNAM9suOGJJZJ4/DJnRIsrjgR8fDhoHcJni4PZCqjAezdc+EdX1Q90LELTnpkXspenauSTTY
pncuT6HIJfCzRCotdJHty38OIOFC+3/EWRbtjrQRqQcytlpn6U7gsPUoObx05hkMNvQbYq6TFSeU
IcH7dehEFrPMLbtHGrA5XmjYvLEIhgQKV9aZ+3U7wUHMjDiof9i6lR8NWEtJAFIRf7Pp6Us2EORu
DzN0N+KAYKuLLb2zOMW3VmxnezDu+dcJv2gnuMyenYVbXrjSSIQAO4Lp8kDwUgd1l1anZut/NJ78
VPnNbLXdkW7VDKwmkLUaX1d2UaFUN67Cvl+q9iM4Gh3H9C3GP25FRSf6YxkPVhjBc38Qm+zO8UJx
5axecRDrR4bBeQsxcZ7KBBcQutbp4rChUJxG+7FlWkeNNYlMZMuNCOLaOdHfQniCOJM4a+sKyVEI
zQvxbXStXQOUoznJDM11gvSbekqQG7wxGKuKFZ+EKA8dMVQnCid138yqSQaAwfwxKGjxtgRnzTW2
G7sBKcb5DGpP1QvBh4qNSy0AeoxpwQsQ+ZuAwuhZiAM2cQHpLwYR1axAWUvjDMzG6WZ5o6VKNUt6
zUTGwe2TayqXNWiPPprytsbN2Ye3uU5uS+1lZCMdVr+yBwmdVqtg1dY+r+PS499vYQi/yqma1W2m
bzn9atVyQBH6cg7Cq9tKU0W9VP1xLVZUoOxBS+WMcO0MTrM8MCKsMq4C1fUbaEO+xmEAvzT3NV6H
noFx6xecHMW8xlMun4kXiQN9Vl8raEbSkQKu0n/Gl5cIHKKeZsasmkH34UyNo/XzmBGrevCwbFsq
NyJANBcalP2ppdBdY6QTHNJ6c9/Kizk6aNKnUC7rRXPx/ivY6tvrHvHHV2hKLCF1Xwno3Fw1hyTk
lrifh8t4lMWx8VKUzhoYW9IW8vrbvF3paohhj/jpT8LTlxRTbgkNRcY49mrtdOyjQx+l0e84J2Mq
tRGPIjSlbP8npHEEORJJGoCi/Cp1NZzHhkdwTW/ezwQAK+Uth2UKNAI8aUkNpzmKwRnXkyxZOvys
PPUPcGnB0qX5R8mVvJT47v94EKVuI4Lt5Ro7flHKrKqge9I1oAZrCgbqQ0whh6yxfXUE5na00ZJO
dhn0b5evcQqsk8WVLASj1xxCyIWdFO9oDP3XcuIwE3WEKxKvwCvHOHNKIyuPpSxcJ0EaccgeEwGn
hdjfXw/C6yS4l6fpK3KqOPX0VHdvlCPUHliC6DPJ1T72IzSNJhMC+lubIl5cyAwEdtLE8w3NUR/G
hYcTCXFJk0aATU8mQT3n0zfhb1537rFJGz+ZsZe5gaNSg62claDsY0ZQ32nB4bh6zgg98xl9oR96
w3Ek8/JdY/R/nUOsp5MYWlLOMCHNR8D0XfP19XA3/cxNy/O3XPkwpgMOvj/Q7R48EnMAUd2LO3Jy
f5g+IwgTAlWb/NbfAKxQZSdCjG7M9rD4ERMYPFncdpJdf7iR6tktyZaa7TX1E2MYXZcinTV2BSiE
9RTts4YIl5680BfAq5R9jE/53Wx61ajmy4+BVRlwXb/FfCPEVNUVvW00MRcgWltFpg71Lk/K0Dx4
pFSrL0r170HYkgAYknENNzrDh6hjrTArzPv/n862/z/YjAlQbW1UcTenZFD5pG3ddQ5AjxYqmhHl
4kv66hZ4sCnctKmRTNjlT2Qsk/mPS60ebrj9TU4uFbYpGj6Ll+Ovd56y2FawYOLnAiLykVBTWL91
QGvlbpbN+hAXKFOiUJQrGpyHQdHDQYx9tMn2yjk94tkn3EfByvZGmof8T5S1LgTPxSrMnk7vA9OJ
3ZCmHojLtgBxYiwUr3ihhZja/JL1qWf8V+W0cWlQk4nRX24CYK4NW82+GlqMnUFfEjyiZ9t5XeW3
P27I7pUgcUiAZ1szWjemAG/FBgmRCjCm/1u+hVqEbn0iS+jcgZu9OGMwhSQaHLBIyF+k6vY1K8ZV
rXTCKyZhxuYvXq3BUSQMrNmmmzAAbiVE49B0JYApq7RbY3Z17LpfHnEUdqVRH3mjHz2Z9bGBkEyV
w7AldqkWkbICisPRh+6k1dHLcHRzS860lMAS7hYMO08Tst50W8ZZMJ0CTIjasA+gcnWvSWEHn3gV
Pypi1BJR+6OnftqbSD/itJT+nh3GLutawcv68XDvHEBkaT3rnei3JOyDFX3KQ4vQMZjS913RIv36
CYYJ7+yKfj67aYDlkR5DLC80lqwqoOrI54Zwfu+fRFxtxNuwGOyWl0jxLGSRBHWrrMuJVOowtM1r
YRzAekgV9x74P06CitrnjfE+fj0+MovMpNT7Lg+d7X/NEHw2FwYOU0jaTatxFwL7GAEkgBnRnGn3
rL2ud1bDfX5uSC/YS/DWd9F42FTKVRAyGZ+Do40mCDOHJwJuRxlofHZ5fo8gs5K6tREdUlG9oT3c
yzDTRgwR2/HiFQ3AjKmEe/oIb/v1qC48VFeulCeVRALPGgaSSMUlVRNRP1sdzKTSEy5sgOlokpGZ
73BADy8rtaevVrFEza11aWNIahKacVPJYn7Blut3oo4uyF/bOZhC5U1z+rrZIG7DNmAYGg9ghE94
4+3AYzmAqmpaL1OXrm7BWxMnj865Mcset5U5BOf8Zkt6XYXAKcdLSVrbVXyAcSwJYP7ULoUZNd42
XWM+FKeQ2n4pbo2nlfeRn2HqLIkKkAbnizqKJoukGpDcEAKEgzd4jSkS2Z72ypLfapcFBLLBPGHR
UEJOcVKhPi0vBGAKZFfw8wnz7Lnv4Hhi1U8ULpZgLSDdR6H4YRyDhkY5uE2exvZmTVnZmnEDPPdJ
jqOswMJOnMORZUhUrQjLPBTeH5APpyGwp4o79/P68926ryFs4Da3WzdPGXsaP2xesMl/KWWuMRNV
RRrMBGQuwIZOifbcsl9gipIs+3I5kjB8JM0AOHG1YalHjaHT6GUSZtacZz8TYrfjllDrNejrKzLd
DjB+l78k80C0jmtcqYAAVy+WJjBscjsDakTwpYrmAhKpu4e0Imv2jd594D2nfz3rvP/dxdLH05mT
vDs2DUM+7/NJdS1dwK5XNqnXg87qjGhIH5nONNozYwrPF70/WEU5o0zvjOG90SkrYtRtjdzTrEiF
K98gTuSqn3D4qTIeGPZqBvmpYTTmQ+TuaKtwGXETaQAdYt01EY8uhBUYyNj06n5KgMSEkLDDZHuH
OHVYZoUz+dHFMMjz3rAQPGMCoUj3KFOzBAsocwS2oT/OzREyAewxEhYc1Ct95EHV57wXkfV3vsKL
kkZGv3minmf7n0Qa3eGeLgKALBHt5i3PBe2fxpmuIpugDse9e4ZHLNRWcBirIP75xc0i3WNyvn0t
XFk1yR6HbjP9tHRDdFiGowNx2NxCpEL/jMs7MFNm57EauLmv/0BplXbFbNghfvruT+2FBU6es5ES
h4gdhWJ+pcoWR/qjBolBH8toy3AT24uZgDWYRgeZ2fANwMGKrb4Vh9ftUI0Zq04GPMsUhDn4Affv
7vGUR3Jl4yQLSXBrPOpS3RE03lifH1qzVNBVEkuMH0n1NF2tndvGKVAUTRaNsotGHXwXoPwFNdrX
QLtvCKFNXP83eqMcRqKUuUdLWdJleXwhTdmYPFV8SXGJOTL4MWiFHBM3OL4NAQKxuLBZEkKsexwq
+sHTdPDCqN7cEVsjyNx/IzA9Kv3f7I8x5ggFRnUHhFYPafcF43QMgtn1mFJBNjqmMbbbzmf6E9p8
RutGbmQf1PjGFFIu0s7vAF5Sg23oRwxNJ2U/2APKOvfDbmKeFDsLFZmLbvoXbItD48iSGadJVmW5
cfhO/MgIA3YUc4JCWLjhDNEFeCp9RViVSc+BfxXCFD+ZSfbmBsfxx+30X/lEzgImtMzC6aseF9Nv
Tp6Rq7ijXIDr7EXeSgvPHQcrYvt2848/YhohpEjvBDO9NoaMr8wBYb8+/i57UNWtREYNyOup87uP
ib9PyrF6CIjlrVH57QkQHSdtLjBHdrVYj0VtEW8ef3poaIMbUJncmT/Jls/BSeDQe1C3J36BydTJ
VBHLkYCK0TqLTNtLZGjyW8yR0nQxqqpmFOaw8esrrBh9bU/r8D5MYiRfF/+Hkzw0QZ8qojaQPzKV
nbNjbO+hs4dXMoYWsbjJBtTzxpaqA1rB5Xfge272q0M1PL8su5TU/OUMgMFMBmR0A8dE/iBmYAzr
K6/S4OqeqIO8YikL7IFvtoCsXVZh0v5DIBogS96ENfUpRMP8Md4eUUInc+UqAkggQSjg4lncQOp0
m2UpVjXdBlCMWVkF5yBgVv22gCjmZNvfgdFVAYTBydINeEzrANi0H4TdQJ3pTW6sgFqsCticLTpN
UOaZBxxMuXopuYbctDONAvOSLxfeK1662RbWKdMKajulPIJUBLw3/ZNS72gUoVKoichehfEgb270
XqL8bgzuSSXwqD/dq314qkKKXIWotMNxo6B5dMK1ltV2vxsQZECWTMd10I656GoU/HRWUUq/GWE6
aSUSXFpxmRBl+Ml5Yb2A2ICa5x60S09itpL0L+xRG6TBdzFiYmIsRuh9VlGXUIx/Bb+r9t9L/S7s
MXeG63QVwXy1qPfkdqHQX4ww8cFuq8ZSgUuDJh3MJPWFH7nbToGX9hprjypvExnDj4txphu0hHF8
ivgBIl8MxXoz2ctP3KgiqC7o9m6oOqPg1K/MZ2AZO+InkfDKk4/iEdMN2ldtuP30+VD9Ae1EByCD
sIL5axTcqP7PbygwbYH5EMGhkLAUOJtR2OoOyaX6/LYcBjynn0fTWl6vgkuYabRf2IEiUFFiW8wh
53q/fRDeUD6VYiXJD4DD3OnPeke/JWAfpcARSyPXwheUkcqLEpJuy/HAgsfL8ErIzQVbcZOVtVPQ
FTgk9FKWZ5buBWezgCW/6zeT9XOZ6grsnV2yPoTdN16WtNF6HpHWZ0QhrylHBnt9qjEtWTjwbZyB
SXFyUvH67P29JQeIzYv9o1ABYS5wBjuSmXIQcM8QTLLWHF3c/wgpG/ZZ5cN/cRmFWzclg2X/alpt
Rpw9rWDnUUYtJvtIjIZrsLY3Sho0odDOhq2PVkP/XAFIBjw+QHH1nb8Ghk687HNEngyzpJaZ8TQm
bvI7TSayLFjtQNLsXqJCSEeCsRhr0Bmwf4FM0+4LbpTvjPmrczFQ1f9rv7b0ypQBBWBdKfx5hlGa
BN3dw1AZQbixXcG7nWnlSYCzPAulcFbOddpADgYrbYYKY6RD7BDbb94Pko6po1BpWKIVYQ6TZH4d
PU+dboJ3E9EU+cKPRW3yaCl+Yn+xrxpdHZJf9Tx5T3/ac2Wd8Sb6dc6y/3kcv400Bkwm+H4KMPhP
C907jOsY1NXB8I68Bs6dHzd+qSKXIbBfRpqGrJVRaD13MxnjCmxizOan3tEID0IztKZVitFs1Iq/
xuOO+teLwsc+FbnNtnxflU5VVtWZRu/Cns8IOaLirwxxKa0ifDtNxCR7Vsdmk60Z7QDO0OUQuk4c
vCYHE4yoU6RZlwC/T3RjPduGmZsXr9mAHa07V1mRrlo9zUTjYRZ1KjmQbLzymCPlHwhjp5YR7vR/
KJk/+78hjgIIY39HgrMtIAjDTN2dseYjNUiNG8hQgVSqFOMmVjrtUqXGNoPdEVyJO36rQeGuAOx7
B+2WZl0uN4bIgPMlmDSks8cUa/wjEWGO8t+n8LH/GazuOjjitk/ZaoQOZFAHB6Giw0hhmB/Tfv8Y
yc9r997sjfIGVvgzsADHAtyvVmQlF3zK/GPkoXqHzfTho8I8rADxURl/y16FlTmqBC5KN+QESF4p
prTroUWdtmZN8KEIBfU5xRRxGhHgb8r3ylYBFTPfPARXEtGLpuaZa7g8x78GbXxSLD6RJoktTX/y
K+87G8QGpdq7fdCHHneqrjBPi7jZXL58HLsoV/wjAuOsUQ/Oif7M4/3w3fw0OJ2FyQ8fV2LCvNyE
LOTt/ukVULxMpvY15vm2aUzlnf7iHbO3ITPIjvCgvxMeUMfjb65GCjzQZ6t9KEmN/9QFSyVaSiKC
9BUi4VUu1ttRUvfq5guW8PrIojLdjiBYvJHY+bAZvBdoOjOzIxh1n2JSx3oZS8P7CHzYz2nNxPGY
G3h89YLG+k0vI51pbF9e/DX2v4cFdQeTNMOW6rFC3mev9TAscxsPhLLGYDKwYyAFkKmfN+SFNcpk
t1ccENm2zamVAxQhei8xZcDpERjARnZsndSFKZ1HZIrKFRuC5LFYXAEYVjpJgG1vAkOb/tMgw5gT
HBcbwNd/o2BC6t9AVVA1hQGsPyfAQnRTUZEfPTB1uNzPUFzacYhPAKJoc4RQG2upfrKMOOxsX8PN
u+My4/G6a133dg4v71BsYFrDEMcJoO5MyaoQzd5VdL1CDEXkO7MaYCada124csN7bCQkX4m6sX/8
Zc5Ld+XxHuaDHGl8woI9zkulIXhJwg+Yk07/WngfHXFP6VKxFclVj+ynFvni976JqfZQsBSugFtC
0XwyNEbXP/TWIcwkj4mZlWRmBqZ2YLeYB+x61cAElV3QdSvuP0eFJH6dcOMuXrBV6kuqztBRzCsp
ueT0N0R8mROxkBEaGv9kG7S6dcTiSEOde/wPm9xbJFcQT7K6S3nqeukQsBxMObhnZZCVmwh4pAJ0
mbUGfpkEKv9TXgNHn5ro7r2vqae+NWU3dYLM8ZhXQUM5P/8MsYaobZ3QNUZrcjfSpfKxaaMgWnyp
LU/yBg+hT1tTIYmo9e2O2CR1LhtppRdiFLNg1vQCkLFofUoZ0LnWAGIduCJBC/59oxyorNFm3suq
g6w5r+peerR6zpUJZYMoY/3H7YC05CHD7Sz8Y7DTJDUOp56+bKDBXl7tO/FBMkd9pO6LbkIZo93V
3Rj4nKTuphqvXTlaVmTangohPLhsJ7EridePLuoUj5WP3sHUcdpwMLJSojDNMcn/FXvH0JEfUO4W
YofU+JBCWF/p4i1PGRYA1yMDftXkkGUhXZWuPY+V2iPAt47nnqvEsSc9dOiOnvApv+Z9HsNkmjlz
611mM/wFZJ4t5Aw5gThh+0gGq/IOucvT+ADXwDpZB5RIB71LtPcZV5wle7oNA2/X1v6nvixo0x/M
l6escWGzNJL9co8h2HgY/BJABso8qBVmxCHve5sEz+hsxCHPBFMoyyr/CE7eIp8GYqQFWboTsAcO
eN8vwZbKeZ7wO4QfumwH7H16sdlBFmNujOioQVicmfDaoxehDW3+9TGIXTbc6YJbfKTacO5z18FW
Fif53/ZObnGCRSNzEGZst3ANcR5l7lU+b24/TMntlB0O19mOmROQCqvm6gGVpoFxEu+fIG8PDjVW
0OVZeLGVuyW/gv96WTqZsHFX12ctaQEYURbCZxiNSpJAgIzDrNjmf3CoTfcWxu4TcBO4Ejfmqajm
eaIGR3wnd8toQzbHhBS9bETww5Xs/Y7UiEpmOp/89MHIdeYZ2FD8mtv/kKLCpntD7QlPgSvCVjKv
PlXz2Yjqca9I3ELTZnw/tnyBu5emRqRNZcOPsi0Cj8mpKX1f79g4tRznpkPW0VfIg1IhOfa1UzYK
DlG68SCIVc+P8bm2CXp8clULRZT4JSbqj9Uf7xfKD3H+Sw33kjmYEQr0ASE7n4rxXDusOvvKVPxp
bPNKnzm5F8GwpeSTGZN68+myyEZL/ZF3u9Lr46a33aI84/pAyB+9uZplBFfMtRdV3D8JpHWQNSOk
HoFcHqdG3Gh2NoGuAH3YGI2kkTr7okdfBXWe/86Hjb9mH5E/XGmisy4gM3wwfdQCl1wSufrekrfl
LM0/5/GBaK+DigYs2I/tsiQw94hFHikKvqP8LNC2M7CnPHMKQINpuFxlxuJHuhPqeSABAnkMw+YR
ACVk+SAs5Tr12ZgXbxyW/uDcL5rK61WstRo5//HsLMTzvt7n4q5uTydiPUz1r7vP1o4LwP+sYP2/
CL3baiq6f2w9Cii1g0LCK2/tdlYdnuVTKPzR4kBurjw0447VNurkSzaCBIJOMJUbvf/2qlii14XY
zXtg2zAo2PVC3UaDNzAC7BJufEHtOQSIV29PE962fehXbW/+F/k77ByFpAcIGPZ3Lh0RrToXth3o
19LhwfWoqbj1ZTCImlQPVukBcvl2bXmVuBWnOX5m8YFdLT2nWQ2ZtLDggKLLdW894gizgrxVOCNj
J0qeTz3QmH6RCM4ViU5lkqCvqFsWb3r8SKZwV8xhWTibzlSbxCHxUinBFiPsFcWVRQdSrAMN/+ZS
tRD2N5VQ7HKMS1sUqPxt1G1DftD89nHdyydy1WidYuOGrfps7fMZ8uRJTNnK4csqr6iJbeRZrN6p
vb9frM1b7RHBc3Os+F67pFPUQ5pAi3CbW+vyT9hU2PD/p6aMO7S+lbUne0CZ8WIZ8zAfsiEQaOmw
ZTyv20gvXasJkTylhpQHC4colz3pvAr9lauISjDQlbEGEFROKmwErsbNHpbrqpEob3+3cPlhcHqX
oEFbmdOqEzAFWjqxnFasd03bfsJmBwG7NynJHmdeieUWOjdFq2ZDg4133Nk7MKQIz1jJuo9E1rtQ
uz5gFfh4MwvPRZedXLZE48eOoX8D37B4wdhAgE0eKboV5AtCh+h0WlAOgCgIvmvidqh4N1bQw6HQ
vi20Ok+oFrjBeo8gMaOi6rUagSnfXNS9d5rByQt9/y1oXnzt6qtcSgfHVwnCBpVAroCfgdxbsXoH
JpQA0sssXYRyKZ/oPPCP3ThtCCSB0IPM0s8+rdSyfEAGkpJwAVro7grBol2Pqb8cOCOkK/08YSc/
yqOJ+A9niaWU52WCRi4h7Xi89AES1xnGN/Zcx4g/pIFcX7KEAqW1ahWTm+Uz4NRbkEiDtEjUJiB4
Ddjfh5/J+5HFs2rNZMmBEG/HDeCUQ3KijVsD37WVfzvhFom3A+aQFZHbHx2p3JECfbDgJGaiM3pk
LjaJJMzMCyIewIwCkCaJKO0v0KG10ubsKaYbojKwNyFjVgtdm9M4BazS4pE4mVEuBNP2PF0SXk6L
gpVEFIRADvR15oQ9TSP/vDK3NEnFE1epKPN359yxYlZP+1umAcsr6oAF+okJEARb7L9L3MxLNqh1
bxWLjhHKX4aNbOeCo1vAe/fQ/crIJsuvr7O4L2nff5UHZIQc5TbpuCLDBVznZUg06aLt0CqqNawc
V2icqZSVVBfKyq9K02FHTVoH0fBwEZdA6dcrtzMhZr0Q8E2get8PM97sha+UawxlbTr01CRuexpv
JwnfZi+179h+YO1B8KLkxCGNktjUxbgR6tiPL9CCJR8Iuasiho/HY3KX9RQWyzMr/TU7vtsAvoZN
g2BHwwVn6RPjOGkuTCg/qudctMtaBu9F5c+5nyuSC91VVsnhn/TLxZ1OuBlHSDfC8vY9xgWJerwM
nvPXy/9AS/69J5NkslY42LuUfkKX3mIXDKSwZaMNbPPmHUfg5kBHr7I39hHYDAozTxpFGBK4q0nb
ni0NgTb0azYGx+N9oyEPn8etW54Kw/uGw8mklMQjxo+pH066yFdI0OoxoLCmgUPel/uwzmdajwOd
nWvNX2LjrqzcjPcTV3T7Qxm5uMSe76c8+A4sHZk8knhaMGOl8O+qW2zAZ3d9GeKbjfhu2vUvddiJ
igIf3jRyDW7yETJaHsg7+q4S788BsBFifzRL7Swa/TCsCk8OPPOjYyAHFBKpeHuGVEcB97FrqmFF
dKj9mnvZmCPqGtbwpU0FSMgxrr2P2+5WjKfp8JneahNI9bSGOd1Q4Ivtp9DG/5xGAYjZS85io/3t
JKFiEKVFyV71p1xct3IrnGuphNfcngStoU+dgg73o3NTBCjrEoK2vKGzx2QoJCOt33+ZOu0OfpT7
52g9C2isbo5WdhRR2enov3TQzQc1Tlgkl5r6BtUvmOMKYZit2bjzY1dLLuujJ/rByPDuBoHQ+UAg
KT3coUkYqLBIPOs2hokEeREuZKe5B/Yg1IaG++02VJOZwHu5z5apjFlz4OcCP81djOF7QgZ3QnuB
F/KVqQJEghN8oGK/F5LnzwwfbCRvpPMQNObtpt00hCAMG1WIaRPFMdHreYsem5me0ZXCa+9z9iS/
oCq2HZkLEmTKOzYcePAmlpn4yhF0X6j6oJvHiV4Cw0BS42mZhTgV6dU4yUV7mmRYPVh1jrtr/4/J
0snunaR70EFiYtdTaz34b+JZIVfgv2ceH473IonkinApKK/RwnoOoI8zlNRpHM6SnNuHV5xdlUzo
ldQGAsSw3xbnXBJrFfAcmviyYYz19Jxx8kDZRLI6rGPdtaaNckQnVUDNq8a0yz6d8ddytwwgbO7x
fbBffRwXbQx7aoKVrYFaQUjZX78cvDT55L/uqsWHMTe0CInt/Q2baibFDoeF2hmZ7Uk7vhuP/kL4
vVDIwwMD/TLIkc63Tc2rm0NS9wlS6FKyDCbRxaYIqYV6a0opz3STy61dGqoSN6WucSPndioIYBO3
RiD99YVAVi8hBiAncvkWqrlc7Gviy2f/zd7m3i7AavJ+AT3AMdhVsHlFcuZzB0lyp3FkwksO5Cnf
Lsxd4Rjvw921PupnsGNWFS6IBD6nd/BmJRRHqpF5iDLX7g0ml7PjEikRnWYSpsiX4UuMagImF4Z8
YGg3RCmlLlDZAynGEq1v7L3L3xpI4a+kE7TkLYvfywNWUYeepuGfsXmXgiXdhAgqp5FjwfqarLSF
vR5m0gK9KLideYN/gnpHNmE4ONd2j8L7tzAUUpyqq/TT2fSdontaumYdleOIX+5umsQMw9VO5ipR
R9STKiC/XYQkuS5QS+DTsBU+yBhHDW1ShzMgv8FT/FvPE0dj+vhTzOo1m/3zQj/bs5NyZPrvLgt3
Sqwh+GoTwkAkQfj9ANTynppX89bcWIcUBjXV4XoiC4plhcf5pjSqlIS0qNtHnatznGM4IwmMdM34
ktcpcEkCH4CJT3Qam/Ean4tADEt15sE+xEmO4dWDkUuCA2tE2SBK/h/aU/PwvK/KlJW6HFqXclGp
oNoUj29h6okmKioqJvNhP9d1ScaKTRrtj0CtrklZBwoox7UeLDMUDoEDAH0zmHg7j4G1YIh+p0Kn
5nIhejitQC0wVX3m2p3XQBijgbgEeLLgju885CXmwH53SH2S7RXomWYezC/vVfB2qY8qUSzRzVEI
aTcLCz4QIyYE/k1DYHssqdVSuzQQVvAVDdAmNLr1whta0IqeVq4ntLIAMizxPdPAKk9qqt4zd6gn
PQliVdVFfZJzsXR6j6+ePExq0aKrbDlDU95xg7wyyCNzgWouBobLBcOBaCQV8USbV3nNriC8nzSA
tED1MCWhBN0oKwjD5XsJqAC6/lE+A01gej0UE6z3fcIFxhS7fjlN/EdBqqfO5ETixZS/oacOcvkX
MkAugasZh8mNJP+uocZDk79e6haEVWMD0ejpcgVcHtm9EPNudkelDEb7vNClhEaViQ8I6boVjYgG
6iXneR+TJ/oTZz/gzIheAX/GXx8bGet4HtyynZOgCxv6lXcBLeQgNUruET2Wd22SPU/cPhY1G2GX
PZ4RkcrpJw+CRkrEbSenya4rVKs43YHy8xPdzMuE+tbwJGbvfI6zAaYSnRxFPrJqAWtWmokfg/Ik
duXTQwcj1xGpDbVrpKVvRzEKXAmmrn4ITDIv7rW68ADBMqCRioEKmPrTakLs7EB4zaCuBxzWCRdb
FhgKWv8mJ/5VWd5mRLsrZrMwkYpsJS4QOdk8uM22eCU1t+JRoDPXZ8kwM3xkzxQsKi8kHn80a/wk
HGjTCiFUe558GcHjfiSXYAfbXIfljgPVRg5u5KHqeUWdlqQe1oQYBnZtvo4D1HwKbGTOhKF/57Ao
g+NlYaXtbL8MYptDHwntz84qYfYxCpSzILl+eLMys5Hjew/KLjdjsNlQuV8Oe/Jw920aWgBPQ2ab
qEYR86MkhtcdGtMHY+NOdKRNxNmYw7Mg6kGkjT7ixHcq1FJhA/OvsiDwxOzhrpTMKRign0z6hdMX
a6yaVr715170SiSfagusWbq375nSt1OCAQ4PyFh2NyjV+NDU7/ojjj85NUzSEmNoa4IF6UTbZlCO
FSwFWjJkF6mZ92WjikqeFUfNmTCJ91fk6BksUxce0+WAtw6NPRcgA0aiLV/0BIYlx/HZXcOxd5kQ
oTG6l+hShTLuRQZ9XBC7fGqquttfWPGZuOFr4GALc94oV4Xxq7fWbWC5lBljsTIOVB8St7Yft4N2
IKtNue06MEJ7u4lBzVa2P1bc8GTUIHzns7Nvv4U9sMNIkC8vLU2iXYtj3v0oao4IczC3Usekn8Sa
ZbT4W6SA8OU3nk/FSLuz5invAQ8yMBzc6qzo1JtzPZjKTAjUHsmC1aB5h92xZlGAfjv5Y9o9yxxV
y7KusiRgdMqgFnb7gyF9/l2iKpeUTC31vGNrKrOQZPd8x10IPzcI5QqCumNsdqD4y00IICCgMXRL
6VjMcV1FW4p9B8jd2ahvmOx4sNZ4w3RwB0bESYFIGxk83CcZS8+XLGp/KWnHKUFacINkDiWIo2CK
WAkHPHzatsj7qozp7G7QzYTbZj7GtZ8dUHSorKzLeL/JQ4rXDhCGJ0tt+pCEUKMYDYp34mwXapGK
m5eGEJWozjP/ibu55phRwk4Gxue1KuWfWlG2P0WCu56nS0U7+IYTvsjhXp3Lwzqj0LNVtK1V5TVH
UIItz3+OckpI7oliKAmvN01V8FAfx9a28xzN1pwrcDMVTsJ/qph4PIDRhI/dGFgcAOqFcBQFv8/X
K8ec74WDCiRBaHzi0bzX46Y5nstPqRiex7KIfyaqKQgQKWy//5ewDzZccFu+TlJlJOZWIrbKAu5B
7zJelCBUCvF2IPFRrFw6iv+ATgXZd9c1g38OSyF2SS9yQLlWGZFvNcsHWgz2Si7lGUaFwKIQGPMZ
wY42qJZB2wMCjDtEQ7dTkvDYA0+6Xq/B3Z4VEHMGpa5RWAJqD/Z8EjNaWGyBsE199xmQIM1jhaLt
ArYgDzUFADkLMDBQOyRjO+u3jPA5/M60BJw05dHIGcx/heN/cIGA13vNTPkdW8GkwcdlX5RvfW9a
cisgBA9pgUTlTvYCiYpXL8gSV47TKVii73XYlOGLX5BOnGaYpBgZKuKxim2kK7/UIC8xsleLZgm7
frESVtUFHGM/IRfGCPdS8I1fFNwaiet4qs3v0/Y46n26BeSpyF1tXMhaZrfLcky+XGTWJ+exw2p1
nJgOBj+eFKak9vX2bum2wjavHA+goqRY3AHrFxvaHzbeuCpgFSMtV6Au3OO9rhGCIxNxLarhSfZz
03s5/o6DemN4XYcxCOsEliVy52WYgrfCzosn5xGr85Bt+6VKsaMOBp08pyRuicQAc37P10D+15qB
8c8oYP6QR7Q94wKo5IiPK9Ra21i9TLe5IMUVuxKko+ZNR6NDFg26iNC7jm6AkGPZfrROrsdyM6Vq
wrB/QMZON1AMIanpDzZEOxB9PLP3VjaXr0XdMk/Zy+29+G5qS9Iwq+qy17Lbs2uypqly+ooWwNJw
2MQx1u8C8jbfPyHQIgorv9bwSiAIfJtw2vF2SguOLlm8aijsIbdYOBKbdwTScX0+1vhpx4CreBOZ
8tMWL+laAItNUx95pdJideQ1Q9uhMFPh68IwsTEHlLVN+ccnhECmYXHQTffuQl4REWhQGw50zlV/
7tMYZEN1ThE3rz/c4yZnjNVKHhABS/DU/EEyMvlRkWTJKD5tVqBSI0CLUbR36JZZOCfwkViNW7nk
+ib6qgjQ+PrdNzjQ/0pcp1WWUjkkjbbeUGljKBXM3+JC1J6CjgItE0B9y6W+VL+G9wNKt0lVv/ei
7Aj244FBCAIeFbrE9eZpJxHnIYxTsBjqqELQBGr4+yX4GT68jlmKfkyZ3XT0223WIk4X2jztf+XH
Hf3J6BblS+AJVzxtP3gYs+0hO7/en2dtZ5Vhjn1yhz8ekNo4gvUZ2ip4BpCmzf5+VxhcmQtmzB48
zLJVKlxqK51WyDqJ1UlosdaUDKJTCJDurcKoMhdrSLdkrcunrnL28f3cU2IghfSkj11/Zkyl3etv
hB8NP5QhN1nt0vgL/dJFnm0GO8YE4YK4ksEszKh5CCGVP/m1QmRh6C2fntvO4BVpdLbVxsmrWdb/
JWD/oA9XBHp72dJDl49OBygJTJqyLcdlFT3awV9mH6RvgNrrFI3iguM3ct6Z08MTQbvzJRRVtT6y
xhrpubS9lIl/xkHwNE36z3SFGmOQ+Aivs1sD0yxSeLTuPXRt3FNqeuQrgS/cvoGU9NUe3JBSMJ3w
ziBjwz6D4hGruo/SaTcXCGz1eLLkKT1QG1wn7wHNlvSwU6EqH7Xdmpd0slt+ki8VTz1d6sSb6zMv
peU6HUbcPygDuPVjpuOcKziY86mjHetDOFk2RCRpbJuiPxvKQGt1IG4S/zteC4WfIEypXdmOHO6C
N8HU/iZiZeTtxQceU34YFicEiRxxOUZzgOCP3GvOiCoVbKBpjcx3DIBw8N3f7XMLF/DxvKqqte7f
WqhWDvX9/FOaukTd5maGSyQMC3V1NHL2uCjEx7Cb7NWHrZ2RT1XYJB5jOWQYX6AciGm1UwodcBeV
c/OPfx8AqC7Hm6FyK85xcqd2OvWHCybyJwy2Ev30rmUYGmM39hkJuHAdEE7MrgPgkOXetS+ZTM1U
49JfN4fk6rEUzqtyShdYh0mpaaX7e3bDYRUrQ9HsXY4rRkQuIfzl5vGmtyT96zvxVl7HqA2JNfNw
5uwFAOTcN1TsyUVM68ojVkE/Lc/JZzZuql5KvclggJvox5K5sqd2Uf4sgvdP2ZmQu1cQQILKdxgr
7eW7khOZ5OYnpGpD5cWUUU3RNv5E1GfbNkgisimM8moMo7sX3CbFSClem4X2oSGEHAxvYt519fhG
y2AFHbcb7JUyC51ypGL/PBgEOQPTZD5Jvqcsm18ooBN5qa9tXMz7m3ep7N4sQPF6BLn5BRJUQuYb
JmmYoRSfvwv9m4GBZjhINEvD+rGruJ4A7MDGEBm/bw76qjT+OHhxlE5twlYt/cgjVXEYrXIzjTOM
8LWPCtzfRJk2GLSMICBeXdN/h9gU7YSIaTZ1iTixWAMnlx5A+OkVpJqWTroPxjhR6iICFoXqsLk5
DcV8s2TsYJDg9r0R7KV2vawSiycxmD46ixBu46FDLTRa/pLiwRQxvo4ZxhN083lRiyultGIqij8y
pOXrrSrj7YMXR+0UD19xawrPTduPqC53XPwlKiZYFkpeuyVqxb3QfZMH3rhhe8ZBmQTjp5mzVpQa
SvbRItnNsypwg3k1Eoj6Ybik59rIt19e9H6uNxy1LNxPSsXNQqMmr9OH3cBpUbzVek82hAOeyYQN
1U10OpqjI5nj+DdGgM5fYSHEFCmCCJGlaRmuaaAvgptsZ8WQPM7doDtxCTyUlQmvd+b9I/zLuDMj
0tSDpL2kI6+Pjjxw9mbJ+/rkcYPJ2FV8yeaOQho22hUSaCgLM2cvO5Xd5NKnBOR7qygn6fmw7dOx
9rSQF3WvwVpHEwSLzHEdq2YpE3Us2Og9ty/TtydvCCFSc05eqpA6wXVFZWD3hCHkiQMrNS4SKI0I
unFF1DpCBASu/92rsA2uA6Sv50gohw7Jix1YSLYB/v+P7Qp1Ex6gEzS05MhSRWqldj9JuZ9j+qG2
OSvS7einoKr4Ke4sNijR/Ypq10tDmNL9pkRtZzw71FDCnKCizQE0CqbGDb01fjQHlN7SsUIsTOij
8swRE477lZ99urPqp3xqkrp9ZMsp25J9KRTqx9cZ92SjW36BnFnulq9tS4OjOfCgtjb4Gw7ZeJhA
EyCHAWC+dfniwCft8N11aX0DloNv3WZja6iFwnzHdZvIsF5mnGLDp5/fvqNTNMoQKIyha9cYP/bT
xDkAQUr8kpFVoZeCwsj0BybD9PVrBnxEEMcRzscqz4cMuDNPIB/T/z/0NgF8zfHAJY61QzPTXP9G
n5rl/Es99zK6LzaWBWuG36NINxyKfWoHqu+I1OsEMnzVGkLohik86EGoHQZsD2aPtcLBQ7bPjUwG
692sTy1gpoHwCAtdXnHh0SY8SH4syXn9EYJPGKT+gInyPYhP41TKdd4M1FctHU+rRMuq69k0BN+c
mnpjOXVKGcJSvPmuuNuX9oXD0W65Z8GvEvH3Jkz86XpaSZLH+T48+RZVi3lXOjdnwLatMdPbhgax
f0y2sIfjBIi69ArjqpTe4dtqiziQ94jt9tadzjUL62Qsq4qmjqHxMtHOqMbDPDEjIjIkeRSt+Eru
47ELmjI/RjRvkAbhwI3v3uUKbe77EqbiR9lGKYg7W1B3h8XYTiDnpV2qdVab3bpT8CwaEZokSZjO
ncOwlPkoDAPGkTujjcPw33u9ilk8lGzRclkAedzXKEv97Hdho5ry6qLc78Q77P1iH8AdnUeAgG7q
P8hynjLq3goau+8J3mofzYBWQTqfKfmZc54zycVC1e4fmQEFmo/WSusK2sxOHLR2TmN56Exvh7on
7r2GgsXRXRnEmNZCY6ZvpbfXd6pJpq6V999fQk7Pg2BUO53Xbwe4ArgD0o1YuPJux0A0SwSPzLB0
hqEckSPd8zIOxYltIgXDA7/s5ddenhk2y7ygL7kAgj/i4opN+1RJVuFcCv8GtoGQLAptXDsxOMUB
EdAEBstV8PV04Wo9L3943VZDL2KPFz55qDW24X+lLVp5Hc4V67VmVKex3m87+9oXAmFMrbGgYV8M
bd0fVkp6NJ+lm6qp9Ok6X6ahRMKkP3yTTLOpFcT8C9iWohKlRWuiMGg4NlwDtM34f5sqI3FwTcGL
DJJv8NNjDWA517G7LRdpwuNfvCa4lySLurVJzyhnvqUq254gEdMawmHP4IfRgM6JoU7WL57z3pIG
lewqAqYglW0KeYDG0L9Q/ScKnNIHvCzhJBr0/LWLCiNjYQ3qGRWXmBrO0kOHik8aBYsEKa7lb+Du
fJbeu8LU1nemKVc6DzDIAh0CFW1WOI/wziYlBR32S5BA0TSRSevOfc01FZ8t6Q7b2wedRRFqAq5h
SdtK6xKO+KNGjiKhPW1Bg5A+YwZ/lzIOTfGOao4VX9ojK0WY+m62SGpbEb9UQ3luAiDQ6t48D9fW
KQkBuC3rYu45C7D0Ibgt1PQTuTxBIIQQGr/4diDHjn7LzztakRQx4XJjFgyvZbf9JBRuEhh6oRjF
fnmKUnz0V0ecxslflyg12Ya3vx0nT4UxwtBJ7gHnkDbUIMThb/ZCAOgNSIGH/kGqYybYZbIBZCTL
TjHU9O3SOVwYoD1F9mn2/ltU1xvrkfZvNT/gYy1ob4YhW1pBCWM5e0dWARvS9Tin5Dfi4n1kRkb6
pNSYQv5v/T5n32XxQ9zcAwlS2bykNkzoblpMFrX4Xcq+I71vLmTCuZ2lcnTQ3FvrRWE2dSWmuK2w
hLDOpJA0/uT+067J8zJs6YtFC9swfoVvIItx8uwJYU1aSlm2dZubgLaaY2i7tZ8tsRvm8FRizFW8
vQw+y8uU054E1MbD7igYPODMSSEJhl0TrpnF0pUcmKtaFUHGWYrjgZ2Vf/M1hL/CDA/onStDNJIp
QVcDB1Yf9a8u0QUNse+X3xbBEI55te4/78JRtnfVt6yu8uAFLBeA7maG0rruPibRGMmRmEgKoMa7
crH2brVLMp5PO6K4NyjxGaq+6P8U4z3/oEIHqCDk3juaZNS3/7vbzpldt0E2I7VyVrFLVmlpxCl2
GlUrqMgxqkVU0vbjbo5ZGpFGSiUHfpCJ85bccNsemZiL3xG7Z7RTHJyEait/CHKqPhYcmI8r+Lsy
scWI9rwwHE1XEbq2nMHB0kKUMTH/IX0c6AyjNujt2fJkmV9o0qN2hOvy7eOCm6vNL0lL2DktLn1I
wa7JIqieCyvvYgAt9gUu0IBzUfSJLjAczU6u5IKQxcXKaV8c9/fuElRqi+I2/fAjbl+D96pARX8m
8HtAPZieZx1lp43q5RILJRNzRZVagWzL1Lrs5knemafFGZYQ2yz3wLqVjMkuXxbWDoHfkR6S0GzI
ju3yjL16dV7pq+UBCby+0pts/h6cwH/fUA+6xEFcfr5NtoRsQYhVQvXZ256wzokkNAfBWItDK9/E
YrXSKJ1uEs34+9zg9+g21RAtVTqRN4rN/wxYcgL/ZmeHZTZSz49cmZcxeNXOKbAYImJ17tN5V3nb
UxxTPXBkxdQLE8tiGgAQJqH4DM49XAfQrSBWhcOLApm8tKxn1RaA+lw4c9jCOd3EYcWMxHKgnaWZ
wg4qt/kLpMQpOvA2C22K8RffRrlrNa/ezpqXIMTvrNY/mmub5+sHTP4d6AjLj+JXpy1vTAJC+CNW
VeLFzWz62JKJI0fAajAk+ZqrCAWOy6DEptFJg2DvYJnduyd2Yqr1X77qytQGDQMbyr2LqBT/vynX
HEaQ0DJLFE+8qWxXVSd7TBZFXimwkaVOYCZtJu1L6j272tmVetSNDzjz/HwF4ZoSp1SMY5/iaiVb
Cy4IDfjbvm3ad4PBdaXnTMA5DNAusnSHg/xmvmv9/L/Bxu/kz6yBjcf86w8/OhIl5zmt779UuwbR
CA8I4NwOpAcsowp/RcEoTowMRv/boGerfsh4DAyCV2SoSeDwq4yKT15eGyJFwl4wC0UgIUucc1Rc
jQXhmmwKcem5yUQiWvcexV+nL9+Nb+J7fPvkBFhCnIK2afhm4nrcGxCASoz0ucJ+nfjCXlSwMueZ
pgz4oAvNlUaaJc+C4r5168JgKMSzqbsGBmKUBs812JQBS8fVvHqRFGgDFwGigp2nyKWWUeX/jD7n
MFOnz27Ue2X0ApV2AM5J7wiy3frsdTP+th/DbvIbFADeuWH4WZVFB5cOSq5H+x9bFiQWlZHuHvVT
qWs2c/8VvupxSVKhEvqGhj/bshzW/mH5GW93UKsw2WMQyQuFgsNIgtJm1tQf/4vbGQF98Mxd9C1O
R/L6ASDiUEvA7tu0kbOL4FutSi0/d+va7Z1vRRwqeJnx2SxtrICz7W6j7a22qfhkrj0b5RAphIvj
wOo4sX5RA8qyhzuMuu22gdTYax3eh0BXCukiP6t6X62qcp+G4bsm0aAgnkl0e5Q/1Z6cS5xVGM62
hLzelOUdx0HHQftsK8fwFWot0sPzIMOLC8O8VeOEA8kzaEgxoTbTD51dKwxAU7w2DEs+1peuGmTZ
xF6cog3fpKV4iLXlZ2Rc04zTDwhSnL/ep1A7GUihokdltdlJduDWRt6YpBZtHfIa/hFFIUcsYwEE
Wpqr5JecDZ2ZDRXXvqzjrWQ3fn2D4c6r0V+32eTuGS5Bil65nVMVNw6Sx6XwPe4SjWR3QSIwvrXv
H6fAX5ZxYchELj3CJoT0+Lym3GWyFR9hsthdbIq+SGWIh2UjBT0u43MNqeHj+eR5eZEiXq/obWLJ
gc9HB18hsAkDXXOaZnstkQskVo3vtZH2IElvtnGdm40cObfraA7KIxHPfnSzfeGP9hHYsezvUj8o
oGfpEri3KyJ7xrx/MRZPIGzl5JaqAQJnYkdOFXbAQ456ic5rsK7YONgtABZWDRgDreh+sFX3Qc2g
nP38YQHXoyrYvhkv0SFHWvbfQ3tC5KPAt7cCynl+MKZo8I1jdzn3cgD/EJmepyJ7juhp1ktQG/PZ
P1/R8VexWQIjA2H+wsUzgyvTy93UPstq2W9cXXdi33dNA4I+sFUDFKsrllxC3OImn68NA44yls8B
WQD+terGxT1DOafpx5sMPwb9orv6opVihb2btoAdDp4xV2tafzzxXNGTCY06W7XEmN0bahQ0AiMv
QHlxBA5IkMrMmKdMD+SIxPaaUQh73MNMPwJ73GeYHzuXIqv/e35gQBS7zwPqeGd+nGtpJ/7ZuASe
HGes/tsON4Dm0ffN1iBSUhfRjHaAsdwND1NdYGvG+Kpnyh6dggMNsphDxmIK2ZDJvIgfQr5Bvhur
BYom2xECTdYD71D8OqWRqWqNE5J6zG7Jvosaai3ETL7HgIxpSAAmA/ehsyMdw8u5qb2Jx9ktL48S
ZrGEISJAJL8FJKGt1iNx7jngUXWjOwiOSaB53v1PZRazTD35eJzG/Ab1LFNpUU2sUMyo4AbinPkV
R0ciNpVpsswVSnYyqgTE5Z8+k+UXzPeG+1Bc0uJt9WJd28qYVe8Cx7BhFFH5ScMdDRTGJMCUGDTd
bedfjrPh9XsX3lIcnRhOE1MZieAkAcKgLpjBh1gIubX8Gk0E5hQPVs3EL7+LXANGUq9H7j3di3Vc
pWl0h2Kc+ylBsmJQne5uIQzfRhDTHbE7XN4zm2MA4FRp+JJJSzUhaBzfiGmd0RcbSxCp+HePHWIT
BqV109gL2o0BEEJKg8JpyxCxKeyPTxaNtGu1jtsSW/PVc6pdGw629KdUlXVWejGbrGCnlwIHn02O
tR4EvPFH1DL1lsDqSNtfhuZ8uodmm/gmNIPQqbh0w0AbQSMfAt/1QH+C/M34pj6LpuKoSHCNzD4b
5gh4Y/T3Q/Qb+7siNqgcj+/L6BcF9FoC0t7no3KskWb9c8wvXkXIzHkjfDIGjcwZ2+HEX4nn163A
eq4COh9LXFCTpteLm+2tOUpWmcG0Bgqla9dV4Sd9G099PYVYQd9/mBK9jSeeHUJ0jtMpDLZtEtH1
kSe7/i5ErJtqojVc8SF7xIv5k/jY+0YSaYykUxz2HBL3aQK49UjMKyJzb2JVeslu0fdNF10N43mU
1PxIML4sk6stMo9GFRJpVwDRljSsQHjBKK1GV3qB5xlH3gtNZ71CkEIRhRq+bbpCL3jtJS6siVA1
pQDbYYtDMl31xfAnQ/AxooFcXc+hvwry1OrDADuGJNDvwvWMIfkWrDgnrgXXrStzUBL5vK9E2yOP
kE2kNiam2ruEr3rGsKk5ovIFWkIpj6NDWCUOpy971Qi3hf1s/iWIhkV5Za8gYWvvey3aoojSDRfy
CSVQgnzRd9RVZNtXXPPHlTT6/LaM/AmTV434REJyZnH6GgLx8sojrqSqp7bHu32h0XLlUOo1ovF3
mazUNa9eNw+Sl16D/N6/fSfSv/X5tlWqXSeqBL633Db06m/D96mbF0ysmh9l9LVTZjDLZJfr8F4V
DIdBBZn466p1co4G56Onb7E17IYHcLgstX5EU2mCg3k7CtK/FQb+YvqnYIp71XRKJAZ5DydnjEqw
kYvTsBCptWKtL2IjvlxNa9qr+txw7ZWjGhOc8cjigP1M2be7Yf6reIKH6JmKfW6ktdYe2xCEQcP5
T97RqYagG7I2IalWtGE9r7tqJ6N/PKHHRx06M2QJrYPll/2w0dFxYXl3jSBzlT/A2cvwNGRpXyzA
471+TjUBekgz388avnmycc/727J40GvIEAcDUG2BLFwIMIyNfooUUl6ntWOf/xkaFu12tuJsr0s8
bRY4MNAxgsAfPJatchsKXlpkTRylxa0AMxyvWUwsB/uVMqU/tm99lJx08FEDl/ru+vJseUYQ39oF
pHU/c5kAvMn5kK81pNXG2I0W+whl07c9rHIMUCoJhxJBR0b/s9xEXiEyKTJ1d0NU6yohQttlLEKu
SzgvoUOvh/q7C2fdD/GbstPSx7FIri07rc8DdWvbwROgTgO1yQ0wRxB4GvwmQAOl5ux4LFzVPRti
qwO1zZ2gyImJJHl5hnN3V6cS3WfaFU4Eq/CrSsoq410r16EV4/Hn4N3v3oEqvfkAw13XoYQ5qzEa
YaHOakmc5h5Kty+awapgivz/hW6TRw6rU+ewoYMlcrNccgsO7MtsRajm6RUT0PJjkuHdFSoefYTV
7GVCmUg4Y27z3kcYZGf/yciQ1CnP659ubxjamjGKBN0aTpUFPrCs7flqqXG2cZxt0vcUeHMJNUL1
G5EQCwMYZFDYqSeYkSSHPLCXb0zBau+19eFyk9VcinP6sH519Qpm435fjP50UKBClydeMVMbRc9P
oMLxUCznCLTCiFOnrTdHh+ynM1WkSijufKoHlgcL7m5MOAOSAn5TvtdbqTV4fWDkowOmjUBHF+89
oaK2GDa5CSbM7YPcusS1MxbB652lbcubE6b4C7WlC1d4Sse0qCHN65ryyK/jslTFf8J60mQ73afY
hUFhB71z7gj/AbDNm4UQCdIL42jcZx+KuXMeebXVOPuYEJn0GtfGrqDgySFn6o8j1CVsor8KxMgf
Zd0pAoM5z1sZbKMtcnjUhu2yxpIR9NXTF8B0dVtxcnzMnfSg9GyHQALgDsQ4MzZFUhankLbNh4cN
hkBddS5DR+KkUThBT5gABdxAQfLXQMmjKxmoJLHTB7iagHd0t9BKtKsmmp/0Ir7MhTBcdF3q0y6o
hAbTJ+m8lpNL6v/9MRYt86O9kG/K0N06y+cU0nkH1T6o1c+RWM9pc8k1/p7xZAMQQcmyJ++xfAy3
+TzNIc+WZMBQaA2ADH2B2VDMsI0VxZQHvRHd/gFqDnT2+3pYwPgmB5gcvkt6IfpdFP357cym5aFk
bXQ0w6qPCy4v7UXVx658DKDpbNk26Yagb53prAO0jH7Wohak+0WoA2yIPUiJiOSCUefgebySq8/u
ldPPd4DGpX7V8T40pAkwrgSGbbAHonxTv/GQNbDHDPZQ2pkX+fyk6QsElzwMjO04+L5lzWAD//Vf
W+6Fe8L6bDIqPTNe0y9vlXV6DyeJJZMtcAEiY8eA5HfPM92JlhT80ar3vo5DDq5T9ZqNLk9pPNRc
tH/7bkJZcoktK8ZNHfppGvt7ZPg9+DKygzTEscncl3K1BWRAyifVc72dKpfVDaf400F8Ql9PzOsz
Bs1Ogyb87HL2N53uUrMsaSc3atyWEF+ob0n6wHz7JthkEzuHdPnfUtjZhGh/ZmzJqx/Dxfg4sAck
NgtCgI15ceEUh/6OL8HWrNetDvgw6Sf8VIh1mKVf8E6XGU15GfKxvsKUTeYj4YT8XoEpIwORtCrV
80jzxhT7QcIWR8Pja1P0dHMs8ya9WQzAv1GDi1rWQUCxXaV3l2/GmPcOXE0KAk/WlcZ1IB/yUnVG
ubMtUCHTxjbuk9aHoK2ArIkpF8IR0xaOA0dcQqsu4LOox28hrLZRh3RQqqsKPL1wMJ2BPg6HPMUY
5MXrr6DnCsVJbfsi4GE6qSP58KKTbWRmDZimf2I5f67pCq/tnHGf8J20wCpLa5IELSNsBlCYJORb
q3Jq+6aTgYr0Uys6NGGJM+dPLp5/ltoNbOiuC8rC+D4GZjv/eOg6KTef4NSr3Rs70MBS9oBx0YLV
o5apgeWojBTvEBaBsLj9l2VumA/tsuij0PdJ/MWbKXn3mwyWAyn+P4YRwXrbXeOzC7+NFTTy1Gms
ViUFbKkJa7XS38SCZk9Mt8N+5cUNHk9prUdtGSpgDToDftNF0YBUW0abmDdqIYYst1I+jjf26hjn
wweJ+jtCZ+GbhgPZddjmB5pILHFOJIW0pXS3ibuQ4dDDfK4+lSpRDHRadD/vT25jD7uEZ90eaDfo
L9NpArSfCNvJQcOVsUkzUg9GZFtj5RVSNTY+2+uYW2qY6CfDoZqrKV1JBXV2cvG8D3MFKeUp01VL
v2FHgruapUmpeDL0qSid2mEW1YQzM0Ab6+JisCe4wDq/oeceJt7qJTOJRjEgLg2FQXBAaH/zXFFp
HLHOctdvDxZHVrEnIpXj816cZU1oOsx6MPAnp8szWDmLpVt6YE2gaa7ydlMBg5NsD9z0fKYnf2oy
Oz6w/XafxkTaYcfCHXp/ZL+hie0zIEmHgL4WibmH1OyQCJ+rSjupxau9izs+NIzlslEnSnKZ0/+Y
BsQCc0j8hfhu47IpbWvqW9x1PDYa8y+cA37MDsAKwqajzLWIFGmc4p7HbmCSzsVl+WuEV1nUpnfb
LsvC+7BthAS9TkBxcamhsexfTfVxG+nQVDwbfejuEjb8sfS0K0osPjhXaxSV1TWgvCUyd+fGqvWd
4sFLT1NnQP7KWWd874t6AEDpgP0STgzZEnQT8MuXzQs0qvgqUtLRybRKZxPuXW9lQ4KSl7fv0bpL
h+M1wgUhLg8ek/AFDd724JgYkmTveBS4xHPI7RzSi91+tSaoYMu4BGpRy1tjk/yYWmfB5xHOTjua
vlTARmPEDFfjlq37neemh/n1fBHPSxQ=
`pragma protect end_protected
